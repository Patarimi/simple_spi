magic
tech sky130B
magscale 1 2
timestamp 1676908156
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 1104 2128 48852 47376
<< metal2 >>
rect 4250 49200 4306 50000
rect 12530 49200 12586 50000
rect 20810 49200 20866 50000
rect 29090 49200 29146 50000
rect 37370 49200 37426 50000
rect 45650 49200 45706 50000
<< obsm2 >>
rect 1582 49144 4194 49314
rect 4362 49144 12474 49314
rect 12642 49144 20754 49314
rect 20922 49144 29034 49314
rect 29202 49144 37314 49314
rect 37482 49144 45594 49314
rect 45762 49144 45980 49314
rect 1582 2139 45980 49144
<< metal3 >>
rect 0 43392 800 43512
rect 0 31016 800 31136
rect 0 18640 800 18760
rect 0 6264 800 6384
<< obsm3 >>
rect 800 43592 35246 47361
rect 880 43312 35246 43592
rect 800 31216 35246 43312
rect 880 30936 35246 31216
rect 800 18840 35246 30936
rect 880 18560 35246 18840
rect 800 6464 35246 18560
rect 880 6184 35246 6464
rect 800 2143 35246 6184
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< labels >>
rlabel metal2 s 12530 49200 12586 50000 6 reg_addr[0]
port 1 nsew signal output
rlabel metal2 s 20810 49200 20866 50000 6 reg_addr[1]
port 2 nsew signal output
rlabel metal2 s 29090 49200 29146 50000 6 reg_addr[2]
port 3 nsew signal output
rlabel metal2 s 37370 49200 37426 50000 6 reg_bus
port 4 nsew signal bidirectional
rlabel metal2 s 45650 49200 45706 50000 6 reg_clk
port 5 nsew signal output
rlabel metal2 s 4250 49200 4306 50000 6 reg_dir
port 6 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 spi_clk
port 7 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 spi_miso
port 8 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 spi_mosi
port 9 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 spi_sel
port 10 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 11 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 11 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 832828
string GDS_FILE /home/mpotereau/DigitalFlowTest/gf_spi_test/openlane/spi_device/runs/23_02_20_16_47/results/signoff/spi_device.magic.gds
string GDS_START 174560
<< end >>

