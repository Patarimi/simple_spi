magic
tech sky130A
magscale 1 2
timestamp 1672930029
<< obsli1 >>
rect 1104 2159 18860 7633
<< obsm1 >>
rect 1104 2128 18860 8288
<< metal2 >>
rect 4710 9200 4766 10000
rect 4802 9200 4858 10000
rect 4894 9200 4950 10000
rect 4986 9200 5042 10000
rect 5078 9200 5134 10000
rect 5170 9200 5226 10000
rect 5262 9200 5318 10000
rect 5354 9200 5410 10000
rect 5446 9200 5502 10000
rect 5538 9200 5594 10000
rect 5630 9200 5686 10000
rect 5722 9200 5778 10000
rect 5814 9200 5870 10000
rect 5906 9200 5962 10000
rect 5998 9200 6054 10000
rect 6090 9200 6146 10000
rect 6182 9200 6238 10000
rect 6274 9200 6330 10000
rect 6366 9200 6422 10000
rect 6458 9200 6514 10000
rect 6550 9200 6606 10000
rect 6642 9200 6698 10000
rect 6734 9200 6790 10000
rect 6826 9200 6882 10000
rect 6918 9200 6974 10000
rect 7010 9200 7066 10000
rect 7102 9200 7158 10000
rect 7194 9200 7250 10000
rect 7286 9200 7342 10000
rect 7378 9200 7434 10000
rect 7470 9200 7526 10000
rect 7562 9200 7618 10000
rect 7654 9200 7710 10000
rect 7746 9200 7802 10000
rect 7838 9200 7894 10000
rect 7930 9200 7986 10000
rect 8022 9200 8078 10000
rect 8114 9200 8170 10000
rect 8206 9200 8262 10000
rect 8298 9200 8354 10000
rect 8390 9200 8446 10000
rect 8482 9200 8538 10000
rect 8574 9200 8630 10000
rect 8666 9200 8722 10000
rect 8758 9200 8814 10000
rect 8850 9200 8906 10000
rect 8942 9200 8998 10000
rect 9034 9200 9090 10000
rect 9126 9200 9182 10000
rect 9218 9200 9274 10000
rect 9310 9200 9366 10000
rect 9402 9200 9458 10000
rect 9494 9200 9550 10000
rect 9586 9200 9642 10000
rect 9678 9200 9734 10000
rect 9770 9200 9826 10000
rect 9862 9200 9918 10000
rect 9954 9200 10010 10000
rect 10046 9200 10102 10000
rect 10138 9200 10194 10000
rect 10230 9200 10286 10000
rect 10322 9200 10378 10000
rect 10414 9200 10470 10000
rect 10506 9200 10562 10000
rect 10598 9200 10654 10000
rect 10690 9200 10746 10000
rect 10782 9200 10838 10000
rect 10874 9200 10930 10000
rect 10966 9200 11022 10000
rect 11058 9200 11114 10000
rect 11150 9200 11206 10000
rect 11242 9200 11298 10000
rect 11334 9200 11390 10000
rect 11426 9200 11482 10000
rect 11518 9200 11574 10000
rect 11610 9200 11666 10000
rect 11702 9200 11758 10000
rect 11794 9200 11850 10000
rect 11886 9200 11942 10000
rect 11978 9200 12034 10000
rect 12070 9200 12126 10000
rect 12162 9200 12218 10000
rect 12254 9200 12310 10000
rect 12346 9200 12402 10000
rect 12438 9200 12494 10000
rect 12530 9200 12586 10000
rect 12622 9200 12678 10000
rect 12714 9200 12770 10000
rect 12806 9200 12862 10000
rect 12898 9200 12954 10000
rect 12990 9200 13046 10000
rect 13082 9200 13138 10000
rect 13174 9200 13230 10000
rect 13266 9200 13322 10000
rect 13358 9200 13414 10000
rect 13450 9200 13506 10000
rect 13542 9200 13598 10000
rect 13634 9200 13690 10000
rect 13726 9200 13782 10000
rect 13818 9200 13874 10000
rect 13910 9200 13966 10000
rect 14002 9200 14058 10000
rect 14094 9200 14150 10000
rect 14186 9200 14242 10000
rect 14278 9200 14334 10000
rect 14370 9200 14426 10000
rect 14462 9200 14518 10000
rect 14554 9200 14610 10000
rect 14646 9200 14702 10000
rect 14738 9200 14794 10000
rect 14830 9200 14886 10000
rect 14922 9200 14978 10000
rect 15014 9200 15070 10000
rect 15106 9200 15162 10000
<< obsm2 >>
rect 1584 9144 4654 9200
rect 15218 9144 18196 9200
rect 1584 2139 18196 9144
<< obsm3 >>
rect 3165 2143 17458 7649
<< metal4 >>
rect 3163 2128 3483 7664
rect 3823 2128 4143 7752
rect 7602 2128 7922 7664
rect 8262 2128 8582 7752
rect 12041 2128 12361 7664
rect 12701 2128 13021 7752
rect 16480 2128 16800 7664
rect 17140 2128 17460 7752
<< metal5 >>
rect 1056 7432 18908 7752
rect 1056 6772 18908 7092
rect 1056 6073 18908 6393
rect 1056 5413 18908 5733
rect 1056 4714 18908 5034
rect 1056 4054 18908 4374
rect 1056 3355 18908 3675
rect 1056 2695 18908 3015
<< labels >>
rlabel metal2 s 4710 9200 4766 10000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 7470 9200 7526 10000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 7746 9200 7802 10000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 8022 9200 8078 10000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 8298 9200 8354 10000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 8574 9200 8630 10000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 8850 9200 8906 10000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 9126 9200 9182 10000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 9402 9200 9458 10000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 9678 9200 9734 10000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 9954 9200 10010 10000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4986 9200 5042 10000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 10230 9200 10286 10000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 10506 9200 10562 10000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 10782 9200 10838 10000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 11058 9200 11114 10000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 11334 9200 11390 10000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 11610 9200 11666 10000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 11886 9200 11942 10000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 12162 9200 12218 10000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 12438 9200 12494 10000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 12714 9200 12770 10000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5262 9200 5318 10000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 12990 9200 13046 10000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 13266 9200 13322 10000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 13542 9200 13598 10000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 13818 9200 13874 10000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 14094 9200 14150 10000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 14370 9200 14426 10000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 14646 9200 14702 10000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 14922 9200 14978 10000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 5538 9200 5594 10000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 5814 9200 5870 10000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 6090 9200 6146 10000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 6366 9200 6422 10000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 6642 9200 6698 10000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 6918 9200 6974 10000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 7194 9200 7250 10000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4802 9200 4858 10000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 7562 9200 7618 10000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 7838 9200 7894 10000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 8114 9200 8170 10000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 8390 9200 8446 10000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 8666 9200 8722 10000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 8942 9200 8998 10000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 9218 9200 9274 10000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 9494 9200 9550 10000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 9770 9200 9826 10000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 10046 9200 10102 10000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 5078 9200 5134 10000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 10322 9200 10378 10000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 10598 9200 10654 10000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 10874 9200 10930 10000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 11150 9200 11206 10000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 11426 9200 11482 10000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 11702 9200 11758 10000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 11978 9200 12034 10000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 12254 9200 12310 10000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 12530 9200 12586 10000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 12806 9200 12862 10000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 5354 9200 5410 10000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 13082 9200 13138 10000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 13358 9200 13414 10000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 13634 9200 13690 10000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 13910 9200 13966 10000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 14186 9200 14242 10000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 14462 9200 14518 10000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 14738 9200 14794 10000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 15014 9200 15070 10000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 5630 9200 5686 10000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 5906 9200 5962 10000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 6182 9200 6238 10000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 6458 9200 6514 10000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 6734 9200 6790 10000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 7010 9200 7066 10000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 7286 9200 7342 10000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4894 9200 4950 10000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 7654 9200 7710 10000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 7930 9200 7986 10000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 8206 9200 8262 10000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 8482 9200 8538 10000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 8758 9200 8814 10000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 9034 9200 9090 10000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 9310 9200 9366 10000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 9586 9200 9642 10000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 9862 9200 9918 10000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 10138 9200 10194 10000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5170 9200 5226 10000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 10414 9200 10470 10000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 10690 9200 10746 10000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 10966 9200 11022 10000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 11242 9200 11298 10000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 11518 9200 11574 10000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 11794 9200 11850 10000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 12070 9200 12126 10000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 12346 9200 12402 10000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 12622 9200 12678 10000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 12898 9200 12954 10000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 5446 9200 5502 10000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 13174 9200 13230 10000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 13450 9200 13506 10000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 13726 9200 13782 10000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 14002 9200 14058 10000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 14278 9200 14334 10000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 14554 9200 14610 10000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 14830 9200 14886 10000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 15106 9200 15162 10000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 5722 9200 5778 10000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 5998 9200 6054 10000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 6274 9200 6330 10000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 6550 9200 6606 10000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 6826 9200 6882 10000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 7102 9200 7158 10000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 7378 9200 7434 10000 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 3163 2128 3483 7664 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 7664 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 7664 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 7664 6 vccd1
port 115 nsew power bidirectional
rlabel metal5 s 1056 2695 18908 3015 6 vccd1
port 115 nsew power bidirectional
rlabel metal5 s 1056 4054 18908 4374 6 vccd1
port 115 nsew power bidirectional
rlabel metal5 s 1056 5413 18908 5733 6 vccd1
port 115 nsew power bidirectional
rlabel metal5 s 1056 6772 18908 7092 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 3823 2128 4143 7752 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 8262 2128 8582 7752 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 12701 2128 13021 7752 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 17140 2128 17460 7752 6 vssd1
port 116 nsew ground bidirectional
rlabel metal5 s 1056 3355 18908 3675 6 vssd1
port 116 nsew ground bidirectional
rlabel metal5 s 1056 4714 18908 5034 6 vssd1
port 116 nsew ground bidirectional
rlabel metal5 s 1056 6073 18908 6393 6 vssd1
port 116 nsew ground bidirectional
rlabel metal5 s 1056 7432 18908 7752 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 405354
string GDS_FILE /home/mpotereau/DigitalFlowTest/gf_spi_test/openlane/spi_wrapper/runs/23_01_05_15_45/results/signoff/spi_wrapper.magic.gds
string GDS_START 152876
<< end >>

