magic
tech sky130A
magscale 1 2
timestamp 1673535444
<< viali >>
rect 1685 15657 1719 15691
rect 4077 15657 4111 15691
rect 5825 15657 5859 15691
rect 8033 15657 8067 15691
rect 10241 15657 10275 15691
rect 12449 15657 12483 15691
rect 14657 15657 14691 15691
rect 16221 15657 16255 15691
rect 1869 15453 1903 15487
rect 4261 15453 4295 15487
rect 6009 15453 6043 15487
rect 8217 15453 8251 15487
rect 10425 15453 10459 15487
rect 12633 15453 12667 15487
rect 14841 15453 14875 15487
rect 16037 15453 16071 15487
rect 2329 15317 2363 15351
rect 10333 6749 10367 6783
rect 12633 6749 12667 6783
rect 12909 6749 12943 6783
rect 10149 6613 10183 6647
rect 13645 6613 13679 6647
rect 9321 6273 9355 6307
rect 9873 6273 9907 6307
rect 10149 6273 10183 6307
rect 11989 6273 12023 6307
rect 13553 6273 13587 6307
rect 11713 6205 11747 6239
rect 13277 6205 13311 6239
rect 9137 6069 9171 6103
rect 10885 6069 10919 6103
rect 12725 6069 12759 6103
rect 14289 6069 14323 6103
rect 10149 5865 10183 5899
rect 11345 5865 11379 5899
rect 12173 5865 12207 5899
rect 12633 5865 12667 5899
rect 13277 5865 13311 5899
rect 14933 5797 14967 5831
rect 9137 5729 9171 5763
rect 12081 5729 12115 5763
rect 14473 5729 14507 5763
rect 15209 5729 15243 5763
rect 15326 5729 15360 5763
rect 15485 5729 15519 5763
rect 9413 5661 9447 5695
rect 11161 5661 11195 5695
rect 12173 5661 12207 5695
rect 12817 5661 12851 5695
rect 13461 5661 13495 5695
rect 14289 5661 14323 5695
rect 10609 5525 10643 5559
rect 11805 5525 11839 5559
rect 16129 5525 16163 5559
rect 9505 5321 9539 5355
rect 11713 5321 11747 5355
rect 12909 5321 12943 5355
rect 13737 5321 13771 5355
rect 11897 5253 11931 5287
rect 8769 5185 8803 5219
rect 12081 5185 12115 5219
rect 12541 5185 12575 5219
rect 13369 5185 13403 5219
rect 13553 5185 13587 5219
rect 14565 5185 14599 5219
rect 8493 5117 8527 5151
rect 12633 5117 12667 5151
rect 16313 5117 16347 5151
rect 12725 4981 12759 5015
rect 8585 4777 8619 4811
rect 11345 4777 11379 4811
rect 11529 4777 11563 4811
rect 12541 4777 12575 4811
rect 15301 4777 15335 4811
rect 8493 4641 8527 4675
rect 10609 4641 10643 4675
rect 8585 4573 8619 4607
rect 9321 4573 9355 4607
rect 9505 4573 9539 4607
rect 10333 4573 10367 4607
rect 10517 4573 10551 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 11621 4573 11655 4607
rect 11713 4573 11747 4607
rect 12357 4573 12391 4607
rect 13369 4573 13403 4607
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 15761 4573 15795 4607
rect 12173 4505 12207 4539
rect 13185 4505 13219 4539
rect 8217 4437 8251 4471
rect 9689 4437 9723 4471
rect 10149 4437 10183 4471
rect 13001 4437 13035 4471
rect 15853 4437 15887 4471
rect 8585 4233 8619 4267
rect 13369 4233 13403 4267
rect 8401 4097 8435 4131
rect 9321 4097 9355 4131
rect 9413 4097 9447 4131
rect 10517 4097 10551 4131
rect 10701 4097 10735 4131
rect 11989 4097 12023 4131
rect 12909 4097 12943 4131
rect 14289 4097 14323 4131
rect 16046 4097 16080 4131
rect 16313 4097 16347 4131
rect 10609 4029 10643 4063
rect 10793 4029 10827 4063
rect 14105 4029 14139 4063
rect 14473 4029 14507 4063
rect 9045 3961 9079 3995
rect 14933 3961 14967 3995
rect 9229 3893 9263 3927
rect 10333 3893 10367 3927
rect 12265 3893 12299 3927
rect 12449 3893 12483 3927
rect 13001 3893 13035 3927
rect 10885 3689 10919 3723
rect 11529 3689 11563 3723
rect 12541 3689 12575 3723
rect 14933 3621 14967 3655
rect 11529 3553 11563 3587
rect 10977 3485 11011 3519
rect 11713 3485 11747 3519
rect 12357 3485 12391 3519
rect 13001 3485 13035 3519
rect 13185 3485 13219 3519
rect 16046 3485 16080 3519
rect 16313 3485 16347 3519
rect 11437 3417 11471 3451
rect 14381 3417 14415 3451
rect 10333 3349 10367 3383
rect 11897 3349 11931 3383
rect 13185 3349 13219 3383
rect 8217 3145 8251 3179
rect 12725 3145 12759 3179
rect 13737 3145 13771 3179
rect 14565 3077 14599 3111
rect 7757 3009 7791 3043
rect 8033 3009 8067 3043
rect 8401 3009 8435 3043
rect 9689 3009 9723 3043
rect 10701 3009 10735 3043
rect 11989 3009 12023 3043
rect 13369 3009 13403 3043
rect 16313 3009 16347 3043
rect 9413 2941 9447 2975
rect 11713 2941 11747 2975
rect 13277 2941 13311 2975
rect 8033 2805 8067 2839
rect 1869 2601 1903 2635
rect 7941 2601 7975 2635
rect 9321 2601 9355 2635
rect 9965 2601 9999 2635
rect 11713 2601 11747 2635
rect 12357 2601 12391 2635
rect 10517 2533 10551 2567
rect 15853 2533 15887 2567
rect 13737 2465 13771 2499
rect 1685 2397 1719 2431
rect 2329 2397 2363 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 6837 2397 6871 2431
rect 7297 2397 7331 2431
rect 8125 2397 8159 2431
rect 8217 2397 8251 2431
rect 9137 2397 9171 2431
rect 9873 2397 9907 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 11897 2397 11931 2431
rect 13470 2397 13504 2431
rect 14565 2397 14599 2431
rect 7941 2329 7975 2363
rect 4813 2261 4847 2295
rect 7481 2261 7515 2295
rect 8401 2261 8435 2295
<< metal1 >>
rect 1104 15802 16836 15824
rect 1104 15750 2916 15802
rect 2968 15750 2980 15802
rect 3032 15750 3044 15802
rect 3096 15750 3108 15802
rect 3160 15750 3172 15802
rect 3224 15750 6849 15802
rect 6901 15750 6913 15802
rect 6965 15750 6977 15802
rect 7029 15750 7041 15802
rect 7093 15750 7105 15802
rect 7157 15750 10782 15802
rect 10834 15750 10846 15802
rect 10898 15750 10910 15802
rect 10962 15750 10974 15802
rect 11026 15750 11038 15802
rect 11090 15750 14715 15802
rect 14767 15750 14779 15802
rect 14831 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 16836 15802
rect 1104 15728 16836 15750
rect 1210 15648 1216 15700
rect 1268 15688 1274 15700
rect 1673 15691 1731 15697
rect 1673 15688 1685 15691
rect 1268 15660 1685 15688
rect 1268 15648 1274 15660
rect 1673 15657 1685 15660
rect 1719 15657 1731 15691
rect 1673 15651 1731 15657
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 3476 15660 4077 15688
rect 3476 15648 3482 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 5810 15688 5816 15700
rect 5771 15660 5816 15688
rect 4065 15651 4123 15657
rect 5810 15648 5816 15660
rect 5868 15648 5874 15700
rect 8018 15688 8024 15700
rect 7979 15660 8024 15688
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 10226 15688 10232 15700
rect 10187 15660 10232 15688
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 12434 15688 12440 15700
rect 12395 15660 12440 15688
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 14458 15648 14464 15700
rect 14516 15688 14522 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14516 15660 14657 15688
rect 14516 15648 14522 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 16209 15691 16267 15697
rect 16209 15657 16221 15691
rect 16255 15688 16267 15691
rect 16666 15688 16672 15700
rect 16255 15660 16672 15688
rect 16255 15657 16267 15660
rect 16209 15651 16267 15657
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 10686 15552 10692 15564
rect 6886 15524 10692 15552
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15484 1915 15487
rect 4246 15484 4252 15496
rect 1903 15456 2360 15484
rect 4207 15456 4252 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 2332 15360 2360 15456
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 5997 15487 6055 15493
rect 5997 15453 6009 15487
rect 6043 15484 6055 15487
rect 6886 15484 6914 15524
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 6043 15456 6914 15484
rect 8205 15487 8263 15493
rect 6043 15453 6055 15456
rect 5997 15447 6055 15453
rect 8205 15453 8217 15487
rect 8251 15484 8263 15487
rect 10134 15484 10140 15496
rect 8251 15456 10140 15484
rect 8251 15453 8263 15456
rect 8205 15447 8263 15453
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15453 10471 15487
rect 10413 15447 10471 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15484 12679 15487
rect 13170 15484 13176 15496
rect 12667 15456 13176 15484
rect 12667 15453 12679 15456
rect 12621 15447 12679 15453
rect 10428 15416 10456 15447
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 14274 15444 14280 15496
rect 14332 15484 14338 15496
rect 14829 15487 14887 15493
rect 14829 15484 14841 15487
rect 14332 15456 14841 15484
rect 14332 15444 14338 15456
rect 14829 15453 14841 15456
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 15252 15456 16037 15484
rect 15252 15444 15258 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 13630 15416 13636 15428
rect 10428 15388 13636 15416
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 2314 15348 2320 15360
rect 2275 15320 2320 15348
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 1104 15258 16995 15280
rect 1104 15206 4882 15258
rect 4934 15206 4946 15258
rect 4998 15206 5010 15258
rect 5062 15206 5074 15258
rect 5126 15206 5138 15258
rect 5190 15206 8815 15258
rect 8867 15206 8879 15258
rect 8931 15206 8943 15258
rect 8995 15206 9007 15258
rect 9059 15206 9071 15258
rect 9123 15206 12748 15258
rect 12800 15206 12812 15258
rect 12864 15206 12876 15258
rect 12928 15206 12940 15258
rect 12992 15206 13004 15258
rect 13056 15206 16681 15258
rect 16733 15206 16745 15258
rect 16797 15206 16809 15258
rect 16861 15206 16873 15258
rect 16925 15206 16937 15258
rect 16989 15206 16995 15258
rect 1104 15184 16995 15206
rect 1104 14714 16836 14736
rect 1104 14662 2916 14714
rect 2968 14662 2980 14714
rect 3032 14662 3044 14714
rect 3096 14662 3108 14714
rect 3160 14662 3172 14714
rect 3224 14662 6849 14714
rect 6901 14662 6913 14714
rect 6965 14662 6977 14714
rect 7029 14662 7041 14714
rect 7093 14662 7105 14714
rect 7157 14662 10782 14714
rect 10834 14662 10846 14714
rect 10898 14662 10910 14714
rect 10962 14662 10974 14714
rect 11026 14662 11038 14714
rect 11090 14662 14715 14714
rect 14767 14662 14779 14714
rect 14831 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 16836 14714
rect 1104 14640 16836 14662
rect 1104 14170 16995 14192
rect 1104 14118 4882 14170
rect 4934 14118 4946 14170
rect 4998 14118 5010 14170
rect 5062 14118 5074 14170
rect 5126 14118 5138 14170
rect 5190 14118 8815 14170
rect 8867 14118 8879 14170
rect 8931 14118 8943 14170
rect 8995 14118 9007 14170
rect 9059 14118 9071 14170
rect 9123 14118 12748 14170
rect 12800 14118 12812 14170
rect 12864 14118 12876 14170
rect 12928 14118 12940 14170
rect 12992 14118 13004 14170
rect 13056 14118 16681 14170
rect 16733 14118 16745 14170
rect 16797 14118 16809 14170
rect 16861 14118 16873 14170
rect 16925 14118 16937 14170
rect 16989 14118 16995 14170
rect 1104 14096 16995 14118
rect 1104 13626 16836 13648
rect 1104 13574 2916 13626
rect 2968 13574 2980 13626
rect 3032 13574 3044 13626
rect 3096 13574 3108 13626
rect 3160 13574 3172 13626
rect 3224 13574 6849 13626
rect 6901 13574 6913 13626
rect 6965 13574 6977 13626
rect 7029 13574 7041 13626
rect 7093 13574 7105 13626
rect 7157 13574 10782 13626
rect 10834 13574 10846 13626
rect 10898 13574 10910 13626
rect 10962 13574 10974 13626
rect 11026 13574 11038 13626
rect 11090 13574 14715 13626
rect 14767 13574 14779 13626
rect 14831 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 16836 13626
rect 1104 13552 16836 13574
rect 1104 13082 16995 13104
rect 1104 13030 4882 13082
rect 4934 13030 4946 13082
rect 4998 13030 5010 13082
rect 5062 13030 5074 13082
rect 5126 13030 5138 13082
rect 5190 13030 8815 13082
rect 8867 13030 8879 13082
rect 8931 13030 8943 13082
rect 8995 13030 9007 13082
rect 9059 13030 9071 13082
rect 9123 13030 12748 13082
rect 12800 13030 12812 13082
rect 12864 13030 12876 13082
rect 12928 13030 12940 13082
rect 12992 13030 13004 13082
rect 13056 13030 16681 13082
rect 16733 13030 16745 13082
rect 16797 13030 16809 13082
rect 16861 13030 16873 13082
rect 16925 13030 16937 13082
rect 16989 13030 16995 13082
rect 1104 13008 16995 13030
rect 1104 12538 16836 12560
rect 1104 12486 2916 12538
rect 2968 12486 2980 12538
rect 3032 12486 3044 12538
rect 3096 12486 3108 12538
rect 3160 12486 3172 12538
rect 3224 12486 6849 12538
rect 6901 12486 6913 12538
rect 6965 12486 6977 12538
rect 7029 12486 7041 12538
rect 7093 12486 7105 12538
rect 7157 12486 10782 12538
rect 10834 12486 10846 12538
rect 10898 12486 10910 12538
rect 10962 12486 10974 12538
rect 11026 12486 11038 12538
rect 11090 12486 14715 12538
rect 14767 12486 14779 12538
rect 14831 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 16836 12538
rect 1104 12464 16836 12486
rect 1104 11994 16995 12016
rect 1104 11942 4882 11994
rect 4934 11942 4946 11994
rect 4998 11942 5010 11994
rect 5062 11942 5074 11994
rect 5126 11942 5138 11994
rect 5190 11942 8815 11994
rect 8867 11942 8879 11994
rect 8931 11942 8943 11994
rect 8995 11942 9007 11994
rect 9059 11942 9071 11994
rect 9123 11942 12748 11994
rect 12800 11942 12812 11994
rect 12864 11942 12876 11994
rect 12928 11942 12940 11994
rect 12992 11942 13004 11994
rect 13056 11942 16681 11994
rect 16733 11942 16745 11994
rect 16797 11942 16809 11994
rect 16861 11942 16873 11994
rect 16925 11942 16937 11994
rect 16989 11942 16995 11994
rect 1104 11920 16995 11942
rect 1104 11450 16836 11472
rect 1104 11398 2916 11450
rect 2968 11398 2980 11450
rect 3032 11398 3044 11450
rect 3096 11398 3108 11450
rect 3160 11398 3172 11450
rect 3224 11398 6849 11450
rect 6901 11398 6913 11450
rect 6965 11398 6977 11450
rect 7029 11398 7041 11450
rect 7093 11398 7105 11450
rect 7157 11398 10782 11450
rect 10834 11398 10846 11450
rect 10898 11398 10910 11450
rect 10962 11398 10974 11450
rect 11026 11398 11038 11450
rect 11090 11398 14715 11450
rect 14767 11398 14779 11450
rect 14831 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 16836 11450
rect 1104 11376 16836 11398
rect 1104 10906 16995 10928
rect 1104 10854 4882 10906
rect 4934 10854 4946 10906
rect 4998 10854 5010 10906
rect 5062 10854 5074 10906
rect 5126 10854 5138 10906
rect 5190 10854 8815 10906
rect 8867 10854 8879 10906
rect 8931 10854 8943 10906
rect 8995 10854 9007 10906
rect 9059 10854 9071 10906
rect 9123 10854 12748 10906
rect 12800 10854 12812 10906
rect 12864 10854 12876 10906
rect 12928 10854 12940 10906
rect 12992 10854 13004 10906
rect 13056 10854 16681 10906
rect 16733 10854 16745 10906
rect 16797 10854 16809 10906
rect 16861 10854 16873 10906
rect 16925 10854 16937 10906
rect 16989 10854 16995 10906
rect 1104 10832 16995 10854
rect 1104 10362 16836 10384
rect 1104 10310 2916 10362
rect 2968 10310 2980 10362
rect 3032 10310 3044 10362
rect 3096 10310 3108 10362
rect 3160 10310 3172 10362
rect 3224 10310 6849 10362
rect 6901 10310 6913 10362
rect 6965 10310 6977 10362
rect 7029 10310 7041 10362
rect 7093 10310 7105 10362
rect 7157 10310 10782 10362
rect 10834 10310 10846 10362
rect 10898 10310 10910 10362
rect 10962 10310 10974 10362
rect 11026 10310 11038 10362
rect 11090 10310 14715 10362
rect 14767 10310 14779 10362
rect 14831 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 16836 10362
rect 1104 10288 16836 10310
rect 1104 9818 16995 9840
rect 1104 9766 4882 9818
rect 4934 9766 4946 9818
rect 4998 9766 5010 9818
rect 5062 9766 5074 9818
rect 5126 9766 5138 9818
rect 5190 9766 8815 9818
rect 8867 9766 8879 9818
rect 8931 9766 8943 9818
rect 8995 9766 9007 9818
rect 9059 9766 9071 9818
rect 9123 9766 12748 9818
rect 12800 9766 12812 9818
rect 12864 9766 12876 9818
rect 12928 9766 12940 9818
rect 12992 9766 13004 9818
rect 13056 9766 16681 9818
rect 16733 9766 16745 9818
rect 16797 9766 16809 9818
rect 16861 9766 16873 9818
rect 16925 9766 16937 9818
rect 16989 9766 16995 9818
rect 1104 9744 16995 9766
rect 1104 9274 16836 9296
rect 1104 9222 2916 9274
rect 2968 9222 2980 9274
rect 3032 9222 3044 9274
rect 3096 9222 3108 9274
rect 3160 9222 3172 9274
rect 3224 9222 6849 9274
rect 6901 9222 6913 9274
rect 6965 9222 6977 9274
rect 7029 9222 7041 9274
rect 7093 9222 7105 9274
rect 7157 9222 10782 9274
rect 10834 9222 10846 9274
rect 10898 9222 10910 9274
rect 10962 9222 10974 9274
rect 11026 9222 11038 9274
rect 11090 9222 14715 9274
rect 14767 9222 14779 9274
rect 14831 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 16836 9274
rect 1104 9200 16836 9222
rect 1104 8730 16995 8752
rect 1104 8678 4882 8730
rect 4934 8678 4946 8730
rect 4998 8678 5010 8730
rect 5062 8678 5074 8730
rect 5126 8678 5138 8730
rect 5190 8678 8815 8730
rect 8867 8678 8879 8730
rect 8931 8678 8943 8730
rect 8995 8678 9007 8730
rect 9059 8678 9071 8730
rect 9123 8678 12748 8730
rect 12800 8678 12812 8730
rect 12864 8678 12876 8730
rect 12928 8678 12940 8730
rect 12992 8678 13004 8730
rect 13056 8678 16681 8730
rect 16733 8678 16745 8730
rect 16797 8678 16809 8730
rect 16861 8678 16873 8730
rect 16925 8678 16937 8730
rect 16989 8678 16995 8730
rect 1104 8656 16995 8678
rect 1104 8186 16836 8208
rect 1104 8134 2916 8186
rect 2968 8134 2980 8186
rect 3032 8134 3044 8186
rect 3096 8134 3108 8186
rect 3160 8134 3172 8186
rect 3224 8134 6849 8186
rect 6901 8134 6913 8186
rect 6965 8134 6977 8186
rect 7029 8134 7041 8186
rect 7093 8134 7105 8186
rect 7157 8134 10782 8186
rect 10834 8134 10846 8186
rect 10898 8134 10910 8186
rect 10962 8134 10974 8186
rect 11026 8134 11038 8186
rect 11090 8134 14715 8186
rect 14767 8134 14779 8186
rect 14831 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 16836 8186
rect 1104 8112 16836 8134
rect 1104 7642 16995 7664
rect 1104 7590 4882 7642
rect 4934 7590 4946 7642
rect 4998 7590 5010 7642
rect 5062 7590 5074 7642
rect 5126 7590 5138 7642
rect 5190 7590 8815 7642
rect 8867 7590 8879 7642
rect 8931 7590 8943 7642
rect 8995 7590 9007 7642
rect 9059 7590 9071 7642
rect 9123 7590 12748 7642
rect 12800 7590 12812 7642
rect 12864 7590 12876 7642
rect 12928 7590 12940 7642
rect 12992 7590 13004 7642
rect 13056 7590 16681 7642
rect 16733 7590 16745 7642
rect 16797 7590 16809 7642
rect 16861 7590 16873 7642
rect 16925 7590 16937 7642
rect 16989 7590 16995 7642
rect 1104 7568 16995 7590
rect 1104 7098 16836 7120
rect 1104 7046 2916 7098
rect 2968 7046 2980 7098
rect 3032 7046 3044 7098
rect 3096 7046 3108 7098
rect 3160 7046 3172 7098
rect 3224 7046 6849 7098
rect 6901 7046 6913 7098
rect 6965 7046 6977 7098
rect 7029 7046 7041 7098
rect 7093 7046 7105 7098
rect 7157 7046 10782 7098
rect 10834 7046 10846 7098
rect 10898 7046 10910 7098
rect 10962 7046 10974 7098
rect 11026 7046 11038 7098
rect 11090 7046 14715 7098
rect 14767 7046 14779 7098
rect 14831 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 16836 7098
rect 1104 7024 16836 7046
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 11238 6780 11244 6792
rect 10367 6752 11244 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 12618 6780 12624 6792
rect 12579 6752 12624 6780
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13722 6780 13728 6792
rect 12943 6752 13728 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 9858 6604 9864 6656
rect 9916 6644 9922 6656
rect 10137 6647 10195 6653
rect 10137 6644 10149 6647
rect 9916 6616 10149 6644
rect 9916 6604 9922 6616
rect 10137 6613 10149 6616
rect 10183 6613 10195 6647
rect 13630 6644 13636 6656
rect 13591 6616 13636 6644
rect 10137 6607 10195 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 1104 6554 16995 6576
rect 1104 6502 4882 6554
rect 4934 6502 4946 6554
rect 4998 6502 5010 6554
rect 5062 6502 5074 6554
rect 5126 6502 5138 6554
rect 5190 6502 8815 6554
rect 8867 6502 8879 6554
rect 8931 6502 8943 6554
rect 8995 6502 9007 6554
rect 9059 6502 9071 6554
rect 9123 6502 12748 6554
rect 12800 6502 12812 6554
rect 12864 6502 12876 6554
rect 12928 6502 12940 6554
rect 12992 6502 13004 6554
rect 13056 6502 16681 6554
rect 16733 6502 16745 6554
rect 16797 6502 16809 6554
rect 16861 6502 16873 6554
rect 16925 6502 16937 6554
rect 16989 6502 16995 6554
rect 1104 6480 16995 6502
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9456 6344 10180 6372
rect 9456 6332 9462 6344
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 9272 6276 9321 6304
rect 9272 6264 9278 6276
rect 9309 6273 9321 6276
rect 9355 6273 9367 6307
rect 9858 6304 9864 6316
rect 9819 6276 9864 6304
rect 9309 6267 9367 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10152 6313 10180 6344
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 10183 6276 11989 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 11977 6273 11989 6276
rect 12023 6304 12035 6307
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 12023 6276 13553 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 13541 6273 13553 6276
rect 13587 6304 13599 6307
rect 13722 6304 13728 6316
rect 13587 6276 13728 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 11330 6196 11336 6248
rect 11388 6236 11394 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11388 6208 11713 6236
rect 11388 6196 11394 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 13262 6236 13268 6248
rect 13223 6208 13268 6236
rect 11701 6199 11759 6205
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 9122 6100 9128 6112
rect 9083 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 10410 6060 10416 6112
rect 10468 6100 10474 6112
rect 10686 6100 10692 6112
rect 10468 6072 10692 6100
rect 10468 6060 10474 6072
rect 10686 6060 10692 6072
rect 10744 6100 10750 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10744 6072 10885 6100
rect 10744 6060 10750 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 12713 6103 12771 6109
rect 12713 6069 12725 6103
rect 12759 6100 12771 6103
rect 13170 6100 13176 6112
rect 12759 6072 13176 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 13170 6060 13176 6072
rect 13228 6100 13234 6112
rect 13538 6100 13544 6112
rect 13228 6072 13544 6100
rect 13228 6060 13234 6072
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 14274 6100 14280 6112
rect 14187 6072 14280 6100
rect 14274 6060 14280 6072
rect 14332 6100 14338 6112
rect 15286 6100 15292 6112
rect 14332 6072 15292 6100
rect 14332 6060 14338 6072
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 1104 6010 16836 6032
rect 1104 5958 2916 6010
rect 2968 5958 2980 6010
rect 3032 5958 3044 6010
rect 3096 5958 3108 6010
rect 3160 5958 3172 6010
rect 3224 5958 6849 6010
rect 6901 5958 6913 6010
rect 6965 5958 6977 6010
rect 7029 5958 7041 6010
rect 7093 5958 7105 6010
rect 7157 5958 10782 6010
rect 10834 5958 10846 6010
rect 10898 5958 10910 6010
rect 10962 5958 10974 6010
rect 11026 5958 11038 6010
rect 11090 5958 14715 6010
rect 14767 5958 14779 6010
rect 14831 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 16836 6010
rect 1104 5936 16836 5958
rect 10134 5896 10140 5908
rect 10095 5868 10140 5896
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 11330 5896 11336 5908
rect 11291 5868 11336 5896
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5865 12219 5899
rect 12618 5896 12624 5908
rect 12579 5868 12624 5896
rect 12161 5859 12219 5865
rect 12176 5828 12204 5859
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 13780 5868 15884 5896
rect 13780 5856 13786 5868
rect 14921 5831 14979 5837
rect 14921 5828 14933 5831
rect 12176 5800 14933 5828
rect 12636 5772 12664 5800
rect 14921 5797 14933 5800
rect 14967 5797 14979 5831
rect 14921 5791 14979 5797
rect 9122 5760 9128 5772
rect 9083 5732 9128 5760
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12342 5760 12348 5772
rect 12115 5732 12348 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12618 5720 12624 5772
rect 12676 5720 12682 5772
rect 13630 5720 13636 5772
rect 13688 5760 13694 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 13688 5732 14473 5760
rect 13688 5720 13694 5732
rect 14461 5729 14473 5732
rect 14507 5729 14519 5763
rect 15194 5760 15200 5772
rect 15155 5732 15200 5760
rect 14461 5723 14519 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15286 5720 15292 5772
rect 15344 5769 15350 5772
rect 15344 5763 15372 5769
rect 15360 5729 15372 5763
rect 15344 5723 15372 5729
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15856 5760 15884 5868
rect 15519 5732 15884 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 15344 5720 15350 5723
rect 9398 5692 9404 5704
rect 9359 5664 9404 5692
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 11146 5692 11152 5704
rect 11107 5664 11152 5692
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 13078 5692 13084 5704
rect 12851 5664 13084 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 12176 5624 12204 5655
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 13446 5692 13452 5704
rect 13407 5664 13452 5692
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13596 5664 14289 5692
rect 13596 5652 13602 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 13170 5624 13176 5636
rect 10612 5596 13176 5624
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 10612 5565 10640 5596
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 2372 5528 10609 5556
rect 2372 5516 2378 5528
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 10597 5519 10655 5525
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 11296 5528 11805 5556
rect 11296 5516 11302 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15344 5528 16129 5556
rect 15344 5516 15350 5528
rect 16117 5525 16129 5528
rect 16163 5525 16175 5559
rect 16117 5519 16175 5525
rect 1104 5466 16995 5488
rect 1104 5414 4882 5466
rect 4934 5414 4946 5466
rect 4998 5414 5010 5466
rect 5062 5414 5074 5466
rect 5126 5414 5138 5466
rect 5190 5414 8815 5466
rect 8867 5414 8879 5466
rect 8931 5414 8943 5466
rect 8995 5414 9007 5466
rect 9059 5414 9071 5466
rect 9123 5414 12748 5466
rect 12800 5414 12812 5466
rect 12864 5414 12876 5466
rect 12928 5414 12940 5466
rect 12992 5414 13004 5466
rect 13056 5414 16681 5466
rect 16733 5414 16745 5466
rect 16797 5414 16809 5466
rect 16861 5414 16873 5466
rect 16925 5414 16937 5466
rect 16989 5414 16995 5466
rect 1104 5392 16995 5414
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 9490 5352 9496 5364
rect 4304 5324 9496 5352
rect 4304 5312 4310 5324
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11701 5355 11759 5361
rect 11701 5352 11713 5355
rect 11204 5324 11713 5352
rect 11204 5312 11210 5324
rect 11701 5321 11713 5324
rect 11747 5321 11759 5355
rect 11701 5315 11759 5321
rect 12897 5355 12955 5361
rect 12897 5321 12909 5355
rect 12943 5352 12955 5355
rect 13078 5352 13084 5364
rect 12943 5324 13084 5352
rect 12943 5321 12955 5324
rect 12897 5315 12955 5321
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 13725 5355 13783 5361
rect 13725 5352 13737 5355
rect 13504 5324 13737 5352
rect 13504 5312 13510 5324
rect 13725 5321 13737 5324
rect 13771 5321 13783 5355
rect 13725 5315 13783 5321
rect 11885 5287 11943 5293
rect 11885 5253 11897 5287
rect 11931 5284 11943 5287
rect 11931 5256 12572 5284
rect 11931 5253 11943 5256
rect 11885 5247 11943 5253
rect 12544 5228 12572 5256
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9398 5216 9404 5228
rect 8803 5188 9404 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5185 12127 5219
rect 12526 5216 12532 5228
rect 12439 5188 12532 5216
rect 12069 5179 12127 5185
rect 8478 5148 8484 5160
rect 8439 5120 8484 5148
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 12084 5148 12112 5179
rect 12526 5176 12532 5188
rect 12584 5216 12590 5228
rect 13357 5219 13415 5225
rect 13357 5216 13369 5219
rect 12584 5188 13369 5216
rect 12584 5176 12590 5188
rect 13357 5185 13369 5188
rect 13403 5185 13415 5219
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13357 5179 13415 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 14550 5216 14556 5228
rect 14511 5188 14556 5216
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 12434 5148 12440 5160
rect 12084 5120 12440 5148
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5148 12679 5151
rect 13722 5148 13728 5160
rect 12667 5120 13728 5148
rect 12667 5117 12679 5120
rect 12621 5111 12679 5117
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 12636 5080 12664 5111
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 16298 5148 16304 5160
rect 16259 5120 16304 5148
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 12400 5052 12664 5080
rect 12400 5040 12406 5052
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 12713 5015 12771 5021
rect 12713 5012 12725 5015
rect 12676 4984 12725 5012
rect 12676 4972 12682 4984
rect 12713 4981 12725 4984
rect 12759 5012 12771 5015
rect 13354 5012 13360 5024
rect 12759 4984 13360 5012
rect 12759 4981 12771 4984
rect 12713 4975 12771 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 1104 4922 16836 4944
rect 1104 4870 2916 4922
rect 2968 4870 2980 4922
rect 3032 4870 3044 4922
rect 3096 4870 3108 4922
rect 3160 4870 3172 4922
rect 3224 4870 6849 4922
rect 6901 4870 6913 4922
rect 6965 4870 6977 4922
rect 7029 4870 7041 4922
rect 7093 4870 7105 4922
rect 7157 4870 10782 4922
rect 10834 4870 10846 4922
rect 10898 4870 10910 4922
rect 10962 4870 10974 4922
rect 11026 4870 11038 4922
rect 11090 4870 14715 4922
rect 14767 4870 14779 4922
rect 14831 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 16836 4922
rect 1104 4848 16836 4870
rect 8570 4808 8576 4820
rect 8531 4780 8576 4808
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 11330 4808 11336 4820
rect 11291 4780 11336 4808
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 11514 4768 11520 4780
rect 11572 4808 11578 4820
rect 12158 4808 12164 4820
rect 11572 4780 12164 4808
rect 11572 4768 11578 4780
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12526 4808 12532 4820
rect 12487 4780 12532 4808
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 15252 4780 15301 4808
rect 15252 4768 15258 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 12434 4740 12440 4752
rect 9416 4712 12440 4740
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 8662 4672 8668 4684
rect 8527 4644 8668 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9416 4672 9444 4712
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 9324 4644 9444 4672
rect 9324 4613 9352 4644
rect 10134 4632 10140 4684
rect 10192 4672 10198 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 10192 4644 10609 4672
rect 10192 4632 10198 4644
rect 10597 4641 10609 4644
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 10704 4644 12480 4672
rect 10704 4616 10732 4644
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 8619 4576 9321 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9309 4573 9321 4576
rect 9355 4573 9367 4607
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9309 4567 9367 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10410 4604 10416 4616
rect 10367 4576 10416 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10520 4536 10548 4567
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 10873 4607 10931 4613
rect 10744 4576 10837 4604
rect 10744 4564 10750 4576
rect 10873 4573 10885 4607
rect 10919 4604 10931 4607
rect 11238 4604 11244 4616
rect 10919 4576 11244 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 11716 4536 11744 4567
rect 11790 4564 11796 4616
rect 11848 4604 11854 4616
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 11848 4576 12357 4604
rect 11848 4564 11854 4576
rect 12345 4573 12357 4576
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12158 4536 12164 4548
rect 10520 4508 11744 4536
rect 12119 4508 12164 4536
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 8386 4468 8392 4480
rect 8251 4440 8392 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9674 4468 9680 4480
rect 9635 4440 9680 4468
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 10134 4468 10140 4480
rect 10095 4440 10140 4468
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 11716 4468 11744 4508
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 12452 4536 12480 4644
rect 12544 4604 12572 4768
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 12544 4576 13369 4604
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 13357 4567 13415 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14516 4576 14565 4604
rect 14516 4564 14522 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 15102 4564 15108 4616
rect 15160 4604 15166 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15160 4576 15761 4604
rect 15160 4564 15166 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 13173 4539 13231 4545
rect 13173 4536 13185 4539
rect 12452 4508 13185 4536
rect 13173 4505 13185 4508
rect 13219 4536 13231 4539
rect 13262 4536 13268 4548
rect 13219 4508 13268 4536
rect 13219 4505 13231 4508
rect 13173 4499 13231 4505
rect 13262 4496 13268 4508
rect 13320 4496 13326 4548
rect 13814 4496 13820 4548
rect 13872 4536 13878 4548
rect 14476 4536 14504 4564
rect 13872 4508 14504 4536
rect 13872 4496 13878 4508
rect 12526 4468 12532 4480
rect 11716 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12676 4440 13001 4468
rect 12676 4428 12682 4440
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 15841 4471 15899 4477
rect 15841 4437 15853 4471
rect 15887 4468 15899 4471
rect 16022 4468 16028 4480
rect 15887 4440 16028 4468
rect 15887 4437 15899 4440
rect 15841 4431 15899 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 1104 4378 16995 4400
rect 1104 4326 4882 4378
rect 4934 4326 4946 4378
rect 4998 4326 5010 4378
rect 5062 4326 5074 4378
rect 5126 4326 5138 4378
rect 5190 4326 8815 4378
rect 8867 4326 8879 4378
rect 8931 4326 8943 4378
rect 8995 4326 9007 4378
rect 9059 4326 9071 4378
rect 9123 4326 12748 4378
rect 12800 4326 12812 4378
rect 12864 4326 12876 4378
rect 12928 4326 12940 4378
rect 12992 4326 13004 4378
rect 13056 4326 16681 4378
rect 16733 4326 16745 4378
rect 16797 4326 16809 4378
rect 16861 4326 16873 4378
rect 16925 4326 16937 4378
rect 16989 4326 16995 4378
rect 1104 4304 16995 4326
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8573 4267 8631 4273
rect 8573 4264 8585 4267
rect 8536 4236 8585 4264
rect 8536 4224 8542 4236
rect 8573 4233 8585 4236
rect 8619 4233 8631 4267
rect 8573 4227 8631 4233
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 13170 4264 13176 4276
rect 12584 4236 13176 4264
rect 12584 4224 12590 4236
rect 13170 4224 13176 4236
rect 13228 4264 13234 4276
rect 13357 4267 13415 4273
rect 13357 4264 13369 4267
rect 13228 4236 13369 4264
rect 13228 4224 13234 4236
rect 13357 4233 13369 4236
rect 13403 4264 13415 4267
rect 13538 4264 13544 4276
rect 13403 4236 13544 4264
rect 13403 4233 13415 4236
rect 13357 4227 13415 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 8386 4128 8392 4140
rect 8347 4100 8392 4128
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9306 4128 9312 4140
rect 8720 4100 9312 4128
rect 8720 4088 8726 4100
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9447 4100 9628 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9214 4060 9220 4072
rect 9048 4032 9220 4060
rect 9048 4001 9076 4032
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9033 3995 9091 4001
rect 9033 3961 9045 3995
rect 9079 3961 9091 3995
rect 9600 3992 9628 4100
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10192 4100 10517 4128
rect 10192 4088 10198 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 11146 4128 11152 4140
rect 10735 4100 11152 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 11146 4088 11152 4100
rect 11204 4128 11210 4140
rect 11790 4128 11796 4140
rect 11204 4100 11796 4128
rect 11204 4088 11210 4100
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11974 4128 11980 4140
rect 11935 4100 11980 4128
rect 11974 4088 11980 4100
rect 12032 4128 12038 4140
rect 12802 4128 12808 4140
rect 12032 4100 12808 4128
rect 12032 4088 12038 4100
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13722 4128 13728 4140
rect 12943 4100 13728 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4128 14335 4131
rect 15286 4128 15292 4140
rect 14323 4100 15292 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16034 4131 16092 4137
rect 16034 4128 16046 4131
rect 15528 4100 16046 4128
rect 15528 4088 15534 4100
rect 16034 4097 16046 4100
rect 16080 4097 16092 4131
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 16034 4091 16092 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 9732 4032 10609 4060
rect 9732 4020 9738 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 10827 4032 14105 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 10686 3992 10692 4004
rect 9600 3964 10692 3992
rect 9033 3955 9091 3961
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 11606 3952 11612 4004
rect 11664 3992 11670 4004
rect 14476 3992 14504 4023
rect 14921 3995 14979 4001
rect 14921 3992 14933 3995
rect 11664 3964 14933 3992
rect 11664 3952 11670 3964
rect 14921 3961 14933 3964
rect 14967 3961 14979 3995
rect 14921 3955 14979 3961
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 9214 3924 9220 3936
rect 8628 3896 9220 3924
rect 8628 3884 8634 3896
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 9732 3896 10333 3924
rect 9732 3884 9738 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 12250 3924 12256 3936
rect 12211 3896 12256 3924
rect 10321 3887 10379 3893
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 12434 3924 12440 3936
rect 12347 3896 12440 3924
rect 12434 3884 12440 3896
rect 12492 3924 12498 3936
rect 12710 3924 12716 3936
rect 12492 3896 12716 3924
rect 12492 3884 12498 3896
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 12860 3896 13001 3924
rect 12860 3884 12866 3896
rect 12989 3893 13001 3896
rect 13035 3924 13047 3927
rect 13354 3924 13360 3936
rect 13035 3896 13360 3924
rect 13035 3893 13047 3896
rect 12989 3887 13047 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 1104 3834 16836 3856
rect 1104 3782 2916 3834
rect 2968 3782 2980 3834
rect 3032 3782 3044 3834
rect 3096 3782 3108 3834
rect 3160 3782 3172 3834
rect 3224 3782 6849 3834
rect 6901 3782 6913 3834
rect 6965 3782 6977 3834
rect 7029 3782 7041 3834
rect 7093 3782 7105 3834
rect 7157 3782 10782 3834
rect 10834 3782 10846 3834
rect 10898 3782 10910 3834
rect 10962 3782 10974 3834
rect 11026 3782 11038 3834
rect 11090 3782 14715 3834
rect 14767 3782 14779 3834
rect 14831 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 16836 3834
rect 1104 3760 16836 3782
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11146 3720 11152 3732
rect 10919 3692 11152 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 11606 3720 11612 3732
rect 11563 3692 11612 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 9306 3612 9312 3664
rect 9364 3652 9370 3664
rect 11532 3652 11560 3683
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12529 3723 12587 3729
rect 12529 3689 12541 3723
rect 12575 3720 12587 3723
rect 14274 3720 14280 3732
rect 12575 3692 14280 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 9364 3624 11560 3652
rect 9364 3612 9370 3624
rect 10980 3525 11008 3624
rect 13354 3612 13360 3664
rect 13412 3652 13418 3664
rect 14921 3655 14979 3661
rect 14921 3652 14933 3655
rect 13412 3624 14933 3652
rect 13412 3612 13418 3624
rect 14921 3621 14933 3624
rect 14967 3652 14979 3655
rect 15102 3652 15108 3664
rect 14967 3624 15108 3652
rect 14967 3621 14979 3624
rect 14921 3615 14979 3621
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 11480 3556 11529 3584
rect 11480 3544 11486 3556
rect 11517 3553 11529 3556
rect 11563 3584 11575 3587
rect 11974 3584 11980 3596
rect 11563 3556 11980 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 10965 3519 11023 3525
rect 10965 3485 10977 3519
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 12250 3516 12256 3528
rect 11747 3488 12256 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 12618 3516 12624 3528
rect 12391 3488 12624 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12768 3488 13001 3516
rect 12768 3476 12774 3488
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 13170 3516 13176 3528
rect 13131 3488 13176 3516
rect 12989 3479 13047 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 16022 3476 16028 3528
rect 16080 3525 16086 3528
rect 16080 3516 16092 3525
rect 16080 3488 16125 3516
rect 16080 3479 16092 3488
rect 16080 3476 16086 3479
rect 16206 3476 16212 3528
rect 16264 3516 16270 3528
rect 16301 3519 16359 3525
rect 16301 3516 16313 3519
rect 16264 3488 16313 3516
rect 16264 3476 16270 3488
rect 16301 3485 16313 3488
rect 16347 3485 16359 3519
rect 16301 3479 16359 3485
rect 9214 3408 9220 3460
rect 9272 3448 9278 3460
rect 11425 3451 11483 3457
rect 11425 3448 11437 3451
rect 9272 3420 11437 3448
rect 9272 3408 9278 3420
rect 11425 3417 11437 3420
rect 11471 3448 11483 3451
rect 11514 3448 11520 3460
rect 11471 3420 11520 3448
rect 11471 3417 11483 3420
rect 11425 3411 11483 3417
rect 11514 3408 11520 3420
rect 11572 3408 11578 3460
rect 14369 3451 14427 3457
rect 14369 3417 14381 3451
rect 14415 3448 14427 3451
rect 14415 3420 15700 3448
rect 14415 3417 14427 3420
rect 14369 3411 14427 3417
rect 10321 3383 10379 3389
rect 10321 3349 10333 3383
rect 10367 3380 10379 3383
rect 10410 3380 10416 3392
rect 10367 3352 10416 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 11882 3380 11888 3392
rect 11843 3352 11888 3380
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 13170 3380 13176 3392
rect 13131 3352 13176 3380
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 15672 3380 15700 3420
rect 16298 3380 16304 3392
rect 15672 3352 16304 3380
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 1104 3290 16995 3312
rect 1104 3238 4882 3290
rect 4934 3238 4946 3290
rect 4998 3238 5010 3290
rect 5062 3238 5074 3290
rect 5126 3238 5138 3290
rect 5190 3238 8815 3290
rect 8867 3238 8879 3290
rect 8931 3238 8943 3290
rect 8995 3238 9007 3290
rect 9059 3238 9071 3290
rect 9123 3238 12748 3290
rect 12800 3238 12812 3290
rect 12864 3238 12876 3290
rect 12928 3238 12940 3290
rect 12992 3238 13004 3290
rect 13056 3238 16681 3290
rect 16733 3238 16745 3290
rect 16797 3238 16809 3290
rect 16861 3238 16873 3290
rect 16925 3238 16937 3290
rect 16989 3238 16995 3290
rect 1104 3216 16995 3238
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 9214 3176 9220 3188
rect 8251 3148 9220 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 12713 3179 12771 3185
rect 12713 3145 12725 3179
rect 12759 3176 12771 3179
rect 13078 3176 13084 3188
rect 12759 3148 13084 3176
rect 12759 3145 12771 3148
rect 12713 3139 12771 3145
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 15470 3176 15476 3188
rect 13771 3148 15476 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 11606 3068 11612 3120
rect 11664 3108 11670 3120
rect 14550 3108 14556 3120
rect 11664 3080 13400 3108
rect 14511 3080 14556 3108
rect 11664 3068 11670 3080
rect 7742 3040 7748 3052
rect 7703 3012 7748 3040
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3040 8079 3043
rect 8202 3040 8208 3052
rect 8067 3012 8208 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8386 3040 8392 3052
rect 8347 3012 8392 3040
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 9674 3040 9680 3052
rect 9635 3012 9680 3040
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 13372 3049 13400 3080
rect 14550 3068 14556 3080
rect 14608 3068 14614 3120
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 10735 3012 11989 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 11977 3009 11989 3012
rect 12023 3040 12035 3043
rect 13357 3043 13415 3049
rect 12023 3012 12388 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 9398 2972 9404 2984
rect 9359 2944 9404 2972
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 11698 2972 11704 2984
rect 11659 2944 11704 2972
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 12360 2904 12388 3012
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 16298 3040 16304 3052
rect 16259 3012 16304 3040
rect 13357 3003 13415 3009
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 13262 2972 13268 2984
rect 13223 2944 13268 2972
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13354 2904 13360 2916
rect 12360 2876 13360 2904
rect 13354 2864 13360 2876
rect 13412 2904 13418 2916
rect 14458 2904 14464 2916
rect 13412 2876 14464 2904
rect 13412 2864 13418 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 8018 2836 8024 2848
rect 7979 2808 8024 2836
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 1104 2746 16836 2768
rect 1104 2694 2916 2746
rect 2968 2694 2980 2746
rect 3032 2694 3044 2746
rect 3096 2694 3108 2746
rect 3160 2694 3172 2746
rect 3224 2694 6849 2746
rect 6901 2694 6913 2746
rect 6965 2694 6977 2746
rect 7029 2694 7041 2746
rect 7093 2694 7105 2746
rect 7157 2694 10782 2746
rect 10834 2694 10846 2746
rect 10898 2694 10910 2746
rect 10962 2694 10974 2746
rect 11026 2694 11038 2746
rect 11090 2694 14715 2746
rect 14767 2694 14779 2746
rect 14831 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 16836 2746
rect 1104 2672 16836 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 1903 2604 7941 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 7929 2601 7941 2604
rect 7975 2632 7987 2635
rect 8386 2632 8392 2644
rect 7975 2604 8392 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9398 2632 9404 2644
rect 9355 2604 9404 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10686 2632 10692 2644
rect 9999 2604 10692 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11698 2632 11704 2644
rect 11659 2604 11704 2632
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 12250 2592 12256 2644
rect 12308 2632 12314 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 12308 2604 12357 2632
rect 12308 2592 12314 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 12345 2595 12403 2601
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2533 10563 2567
rect 10505 2527 10563 2533
rect 15841 2567 15899 2573
rect 15841 2533 15853 2567
rect 15887 2564 15899 2567
rect 16206 2564 16212 2576
rect 15887 2536 16212 2564
rect 15887 2533 15899 2536
rect 15841 2527 15899 2533
rect 10520 2496 10548 2527
rect 8312 2468 10548 2496
rect 13725 2499 13783 2505
rect 1578 2388 1584 2440
rect 1636 2428 1642 2440
rect 1673 2431 1731 2437
rect 1673 2428 1685 2431
rect 1636 2400 1685 2428
rect 1636 2388 1642 2400
rect 1673 2397 1685 2400
rect 1719 2428 1731 2431
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 1719 2400 2329 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2428 4675 2431
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 4663 2400 5273 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 6871 2400 7297 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 7285 2397 7297 2400
rect 7331 2428 7343 2431
rect 7466 2428 7472 2440
rect 7331 2400 7472 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8018 2388 8024 2440
rect 8076 2428 8082 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 8076 2400 8125 2428
rect 8076 2388 8082 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 7742 2360 7748 2372
rect 4816 2332 7748 2360
rect 4816 2301 4844 2332
rect 7742 2320 7748 2332
rect 7800 2360 7806 2372
rect 7929 2363 7987 2369
rect 7929 2360 7941 2363
rect 7800 2332 7941 2360
rect 7800 2320 7806 2332
rect 7929 2329 7941 2332
rect 7975 2329 7987 2363
rect 7929 2323 7987 2329
rect 4801 2295 4859 2301
rect 4801 2261 4813 2295
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 7469 2295 7527 2301
rect 7469 2261 7481 2295
rect 7515 2292 7527 2295
rect 8128 2292 8156 2391
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 8312 2428 8340 2468
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 15856 2496 15884 2527
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 13771 2468 15884 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8260 2400 8353 2428
rect 8404 2400 9137 2428
rect 8260 2388 8266 2400
rect 8404 2301 8432 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 7515 2264 8156 2292
rect 8389 2295 8447 2301
rect 7515 2261 7527 2264
rect 7469 2255 7527 2261
rect 8389 2261 8401 2295
rect 8435 2261 8447 2295
rect 9876 2292 9904 2391
rect 10060 2360 10088 2391
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10468 2400 10701 2428
rect 10468 2388 10474 2400
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 11882 2428 11888 2440
rect 11843 2400 11888 2428
rect 10689 2391 10747 2397
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13458 2431 13516 2437
rect 13458 2428 13470 2431
rect 13228 2400 13470 2428
rect 13228 2388 13234 2400
rect 13458 2397 13470 2400
rect 13504 2397 13516 2431
rect 14550 2428 14556 2440
rect 14511 2400 14556 2428
rect 13458 2391 13516 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 11422 2360 11428 2372
rect 10060 2332 11428 2360
rect 11422 2320 11428 2332
rect 11480 2320 11486 2372
rect 12250 2292 12256 2304
rect 9876 2264 12256 2292
rect 8389 2255 8447 2261
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 1104 2202 16995 2224
rect 1104 2150 4882 2202
rect 4934 2150 4946 2202
rect 4998 2150 5010 2202
rect 5062 2150 5074 2202
rect 5126 2150 5138 2202
rect 5190 2150 8815 2202
rect 8867 2150 8879 2202
rect 8931 2150 8943 2202
rect 8995 2150 9007 2202
rect 9059 2150 9071 2202
rect 9123 2150 12748 2202
rect 12800 2150 12812 2202
rect 12864 2150 12876 2202
rect 12928 2150 12940 2202
rect 12992 2150 13004 2202
rect 13056 2150 16681 2202
rect 16733 2150 16745 2202
rect 16797 2150 16809 2202
rect 16861 2150 16873 2202
rect 16925 2150 16937 2202
rect 16989 2150 16995 2202
rect 1104 2128 16995 2150
<< via1 >>
rect 2916 15750 2968 15802
rect 2980 15750 3032 15802
rect 3044 15750 3096 15802
rect 3108 15750 3160 15802
rect 3172 15750 3224 15802
rect 6849 15750 6901 15802
rect 6913 15750 6965 15802
rect 6977 15750 7029 15802
rect 7041 15750 7093 15802
rect 7105 15750 7157 15802
rect 10782 15750 10834 15802
rect 10846 15750 10898 15802
rect 10910 15750 10962 15802
rect 10974 15750 11026 15802
rect 11038 15750 11090 15802
rect 14715 15750 14767 15802
rect 14779 15750 14831 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 1216 15648 1268 15700
rect 3424 15648 3476 15700
rect 5816 15691 5868 15700
rect 5816 15657 5825 15691
rect 5825 15657 5859 15691
rect 5859 15657 5868 15691
rect 5816 15648 5868 15657
rect 8024 15691 8076 15700
rect 8024 15657 8033 15691
rect 8033 15657 8067 15691
rect 8067 15657 8076 15691
rect 8024 15648 8076 15657
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12440 15648 12492 15657
rect 14464 15648 14516 15700
rect 16672 15648 16724 15700
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 10692 15512 10744 15564
rect 10140 15444 10192 15496
rect 13176 15444 13228 15496
rect 14280 15444 14332 15496
rect 15200 15444 15252 15496
rect 13636 15376 13688 15428
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 4882 15206 4934 15258
rect 4946 15206 4998 15258
rect 5010 15206 5062 15258
rect 5074 15206 5126 15258
rect 5138 15206 5190 15258
rect 8815 15206 8867 15258
rect 8879 15206 8931 15258
rect 8943 15206 8995 15258
rect 9007 15206 9059 15258
rect 9071 15206 9123 15258
rect 12748 15206 12800 15258
rect 12812 15206 12864 15258
rect 12876 15206 12928 15258
rect 12940 15206 12992 15258
rect 13004 15206 13056 15258
rect 16681 15206 16733 15258
rect 16745 15206 16797 15258
rect 16809 15206 16861 15258
rect 16873 15206 16925 15258
rect 16937 15206 16989 15258
rect 2916 14662 2968 14714
rect 2980 14662 3032 14714
rect 3044 14662 3096 14714
rect 3108 14662 3160 14714
rect 3172 14662 3224 14714
rect 6849 14662 6901 14714
rect 6913 14662 6965 14714
rect 6977 14662 7029 14714
rect 7041 14662 7093 14714
rect 7105 14662 7157 14714
rect 10782 14662 10834 14714
rect 10846 14662 10898 14714
rect 10910 14662 10962 14714
rect 10974 14662 11026 14714
rect 11038 14662 11090 14714
rect 14715 14662 14767 14714
rect 14779 14662 14831 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 4882 14118 4934 14170
rect 4946 14118 4998 14170
rect 5010 14118 5062 14170
rect 5074 14118 5126 14170
rect 5138 14118 5190 14170
rect 8815 14118 8867 14170
rect 8879 14118 8931 14170
rect 8943 14118 8995 14170
rect 9007 14118 9059 14170
rect 9071 14118 9123 14170
rect 12748 14118 12800 14170
rect 12812 14118 12864 14170
rect 12876 14118 12928 14170
rect 12940 14118 12992 14170
rect 13004 14118 13056 14170
rect 16681 14118 16733 14170
rect 16745 14118 16797 14170
rect 16809 14118 16861 14170
rect 16873 14118 16925 14170
rect 16937 14118 16989 14170
rect 2916 13574 2968 13626
rect 2980 13574 3032 13626
rect 3044 13574 3096 13626
rect 3108 13574 3160 13626
rect 3172 13574 3224 13626
rect 6849 13574 6901 13626
rect 6913 13574 6965 13626
rect 6977 13574 7029 13626
rect 7041 13574 7093 13626
rect 7105 13574 7157 13626
rect 10782 13574 10834 13626
rect 10846 13574 10898 13626
rect 10910 13574 10962 13626
rect 10974 13574 11026 13626
rect 11038 13574 11090 13626
rect 14715 13574 14767 13626
rect 14779 13574 14831 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 4882 13030 4934 13082
rect 4946 13030 4998 13082
rect 5010 13030 5062 13082
rect 5074 13030 5126 13082
rect 5138 13030 5190 13082
rect 8815 13030 8867 13082
rect 8879 13030 8931 13082
rect 8943 13030 8995 13082
rect 9007 13030 9059 13082
rect 9071 13030 9123 13082
rect 12748 13030 12800 13082
rect 12812 13030 12864 13082
rect 12876 13030 12928 13082
rect 12940 13030 12992 13082
rect 13004 13030 13056 13082
rect 16681 13030 16733 13082
rect 16745 13030 16797 13082
rect 16809 13030 16861 13082
rect 16873 13030 16925 13082
rect 16937 13030 16989 13082
rect 2916 12486 2968 12538
rect 2980 12486 3032 12538
rect 3044 12486 3096 12538
rect 3108 12486 3160 12538
rect 3172 12486 3224 12538
rect 6849 12486 6901 12538
rect 6913 12486 6965 12538
rect 6977 12486 7029 12538
rect 7041 12486 7093 12538
rect 7105 12486 7157 12538
rect 10782 12486 10834 12538
rect 10846 12486 10898 12538
rect 10910 12486 10962 12538
rect 10974 12486 11026 12538
rect 11038 12486 11090 12538
rect 14715 12486 14767 12538
rect 14779 12486 14831 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 4882 11942 4934 11994
rect 4946 11942 4998 11994
rect 5010 11942 5062 11994
rect 5074 11942 5126 11994
rect 5138 11942 5190 11994
rect 8815 11942 8867 11994
rect 8879 11942 8931 11994
rect 8943 11942 8995 11994
rect 9007 11942 9059 11994
rect 9071 11942 9123 11994
rect 12748 11942 12800 11994
rect 12812 11942 12864 11994
rect 12876 11942 12928 11994
rect 12940 11942 12992 11994
rect 13004 11942 13056 11994
rect 16681 11942 16733 11994
rect 16745 11942 16797 11994
rect 16809 11942 16861 11994
rect 16873 11942 16925 11994
rect 16937 11942 16989 11994
rect 2916 11398 2968 11450
rect 2980 11398 3032 11450
rect 3044 11398 3096 11450
rect 3108 11398 3160 11450
rect 3172 11398 3224 11450
rect 6849 11398 6901 11450
rect 6913 11398 6965 11450
rect 6977 11398 7029 11450
rect 7041 11398 7093 11450
rect 7105 11398 7157 11450
rect 10782 11398 10834 11450
rect 10846 11398 10898 11450
rect 10910 11398 10962 11450
rect 10974 11398 11026 11450
rect 11038 11398 11090 11450
rect 14715 11398 14767 11450
rect 14779 11398 14831 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 4882 10854 4934 10906
rect 4946 10854 4998 10906
rect 5010 10854 5062 10906
rect 5074 10854 5126 10906
rect 5138 10854 5190 10906
rect 8815 10854 8867 10906
rect 8879 10854 8931 10906
rect 8943 10854 8995 10906
rect 9007 10854 9059 10906
rect 9071 10854 9123 10906
rect 12748 10854 12800 10906
rect 12812 10854 12864 10906
rect 12876 10854 12928 10906
rect 12940 10854 12992 10906
rect 13004 10854 13056 10906
rect 16681 10854 16733 10906
rect 16745 10854 16797 10906
rect 16809 10854 16861 10906
rect 16873 10854 16925 10906
rect 16937 10854 16989 10906
rect 2916 10310 2968 10362
rect 2980 10310 3032 10362
rect 3044 10310 3096 10362
rect 3108 10310 3160 10362
rect 3172 10310 3224 10362
rect 6849 10310 6901 10362
rect 6913 10310 6965 10362
rect 6977 10310 7029 10362
rect 7041 10310 7093 10362
rect 7105 10310 7157 10362
rect 10782 10310 10834 10362
rect 10846 10310 10898 10362
rect 10910 10310 10962 10362
rect 10974 10310 11026 10362
rect 11038 10310 11090 10362
rect 14715 10310 14767 10362
rect 14779 10310 14831 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 4882 9766 4934 9818
rect 4946 9766 4998 9818
rect 5010 9766 5062 9818
rect 5074 9766 5126 9818
rect 5138 9766 5190 9818
rect 8815 9766 8867 9818
rect 8879 9766 8931 9818
rect 8943 9766 8995 9818
rect 9007 9766 9059 9818
rect 9071 9766 9123 9818
rect 12748 9766 12800 9818
rect 12812 9766 12864 9818
rect 12876 9766 12928 9818
rect 12940 9766 12992 9818
rect 13004 9766 13056 9818
rect 16681 9766 16733 9818
rect 16745 9766 16797 9818
rect 16809 9766 16861 9818
rect 16873 9766 16925 9818
rect 16937 9766 16989 9818
rect 2916 9222 2968 9274
rect 2980 9222 3032 9274
rect 3044 9222 3096 9274
rect 3108 9222 3160 9274
rect 3172 9222 3224 9274
rect 6849 9222 6901 9274
rect 6913 9222 6965 9274
rect 6977 9222 7029 9274
rect 7041 9222 7093 9274
rect 7105 9222 7157 9274
rect 10782 9222 10834 9274
rect 10846 9222 10898 9274
rect 10910 9222 10962 9274
rect 10974 9222 11026 9274
rect 11038 9222 11090 9274
rect 14715 9222 14767 9274
rect 14779 9222 14831 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 4882 8678 4934 8730
rect 4946 8678 4998 8730
rect 5010 8678 5062 8730
rect 5074 8678 5126 8730
rect 5138 8678 5190 8730
rect 8815 8678 8867 8730
rect 8879 8678 8931 8730
rect 8943 8678 8995 8730
rect 9007 8678 9059 8730
rect 9071 8678 9123 8730
rect 12748 8678 12800 8730
rect 12812 8678 12864 8730
rect 12876 8678 12928 8730
rect 12940 8678 12992 8730
rect 13004 8678 13056 8730
rect 16681 8678 16733 8730
rect 16745 8678 16797 8730
rect 16809 8678 16861 8730
rect 16873 8678 16925 8730
rect 16937 8678 16989 8730
rect 2916 8134 2968 8186
rect 2980 8134 3032 8186
rect 3044 8134 3096 8186
rect 3108 8134 3160 8186
rect 3172 8134 3224 8186
rect 6849 8134 6901 8186
rect 6913 8134 6965 8186
rect 6977 8134 7029 8186
rect 7041 8134 7093 8186
rect 7105 8134 7157 8186
rect 10782 8134 10834 8186
rect 10846 8134 10898 8186
rect 10910 8134 10962 8186
rect 10974 8134 11026 8186
rect 11038 8134 11090 8186
rect 14715 8134 14767 8186
rect 14779 8134 14831 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 4882 7590 4934 7642
rect 4946 7590 4998 7642
rect 5010 7590 5062 7642
rect 5074 7590 5126 7642
rect 5138 7590 5190 7642
rect 8815 7590 8867 7642
rect 8879 7590 8931 7642
rect 8943 7590 8995 7642
rect 9007 7590 9059 7642
rect 9071 7590 9123 7642
rect 12748 7590 12800 7642
rect 12812 7590 12864 7642
rect 12876 7590 12928 7642
rect 12940 7590 12992 7642
rect 13004 7590 13056 7642
rect 16681 7590 16733 7642
rect 16745 7590 16797 7642
rect 16809 7590 16861 7642
rect 16873 7590 16925 7642
rect 16937 7590 16989 7642
rect 2916 7046 2968 7098
rect 2980 7046 3032 7098
rect 3044 7046 3096 7098
rect 3108 7046 3160 7098
rect 3172 7046 3224 7098
rect 6849 7046 6901 7098
rect 6913 7046 6965 7098
rect 6977 7046 7029 7098
rect 7041 7046 7093 7098
rect 7105 7046 7157 7098
rect 10782 7046 10834 7098
rect 10846 7046 10898 7098
rect 10910 7046 10962 7098
rect 10974 7046 11026 7098
rect 11038 7046 11090 7098
rect 14715 7046 14767 7098
rect 14779 7046 14831 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 11244 6740 11296 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13728 6740 13780 6792
rect 9864 6604 9916 6656
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 4882 6502 4934 6554
rect 4946 6502 4998 6554
rect 5010 6502 5062 6554
rect 5074 6502 5126 6554
rect 5138 6502 5190 6554
rect 8815 6502 8867 6554
rect 8879 6502 8931 6554
rect 8943 6502 8995 6554
rect 9007 6502 9059 6554
rect 9071 6502 9123 6554
rect 12748 6502 12800 6554
rect 12812 6502 12864 6554
rect 12876 6502 12928 6554
rect 12940 6502 12992 6554
rect 13004 6502 13056 6554
rect 16681 6502 16733 6554
rect 16745 6502 16797 6554
rect 16809 6502 16861 6554
rect 16873 6502 16925 6554
rect 16937 6502 16989 6554
rect 9404 6332 9456 6384
rect 9220 6264 9272 6316
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 13728 6264 13780 6316
rect 11336 6196 11388 6248
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 10416 6060 10468 6112
rect 10692 6060 10744 6112
rect 13176 6060 13228 6112
rect 13544 6060 13596 6112
rect 14280 6103 14332 6112
rect 14280 6069 14289 6103
rect 14289 6069 14323 6103
rect 14323 6069 14332 6103
rect 14280 6060 14332 6069
rect 15292 6060 15344 6112
rect 2916 5958 2968 6010
rect 2980 5958 3032 6010
rect 3044 5958 3096 6010
rect 3108 5958 3160 6010
rect 3172 5958 3224 6010
rect 6849 5958 6901 6010
rect 6913 5958 6965 6010
rect 6977 5958 7029 6010
rect 7041 5958 7093 6010
rect 7105 5958 7157 6010
rect 10782 5958 10834 6010
rect 10846 5958 10898 6010
rect 10910 5958 10962 6010
rect 10974 5958 11026 6010
rect 11038 5958 11090 6010
rect 14715 5958 14767 6010
rect 14779 5958 14831 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 11336 5899 11388 5908
rect 11336 5865 11345 5899
rect 11345 5865 11379 5899
rect 11379 5865 11388 5899
rect 11336 5856 11388 5865
rect 12624 5899 12676 5908
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 13728 5856 13780 5908
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 12348 5720 12400 5772
rect 12624 5720 12676 5772
rect 13636 5720 13688 5772
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 15292 5763 15344 5772
rect 15292 5729 15326 5763
rect 15326 5729 15344 5763
rect 15292 5720 15344 5729
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 13084 5652 13136 5704
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 13544 5652 13596 5704
rect 2320 5516 2372 5568
rect 13176 5584 13228 5636
rect 11244 5516 11296 5568
rect 15292 5516 15344 5568
rect 4882 5414 4934 5466
rect 4946 5414 4998 5466
rect 5010 5414 5062 5466
rect 5074 5414 5126 5466
rect 5138 5414 5190 5466
rect 8815 5414 8867 5466
rect 8879 5414 8931 5466
rect 8943 5414 8995 5466
rect 9007 5414 9059 5466
rect 9071 5414 9123 5466
rect 12748 5414 12800 5466
rect 12812 5414 12864 5466
rect 12876 5414 12928 5466
rect 12940 5414 12992 5466
rect 13004 5414 13056 5466
rect 16681 5414 16733 5466
rect 16745 5414 16797 5466
rect 16809 5414 16861 5466
rect 16873 5414 16925 5466
rect 16937 5414 16989 5466
rect 4252 5312 4304 5364
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 11152 5312 11204 5364
rect 13084 5312 13136 5364
rect 13452 5312 13504 5364
rect 9404 5176 9456 5228
rect 12532 5219 12584 5228
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 12440 5108 12492 5160
rect 12348 5040 12400 5092
rect 13728 5108 13780 5160
rect 16304 5151 16356 5160
rect 16304 5117 16313 5151
rect 16313 5117 16347 5151
rect 16347 5117 16356 5151
rect 16304 5108 16356 5117
rect 12624 4972 12676 5024
rect 13360 4972 13412 5024
rect 2916 4870 2968 4922
rect 2980 4870 3032 4922
rect 3044 4870 3096 4922
rect 3108 4870 3160 4922
rect 3172 4870 3224 4922
rect 6849 4870 6901 4922
rect 6913 4870 6965 4922
rect 6977 4870 7029 4922
rect 7041 4870 7093 4922
rect 7105 4870 7157 4922
rect 10782 4870 10834 4922
rect 10846 4870 10898 4922
rect 10910 4870 10962 4922
rect 10974 4870 11026 4922
rect 11038 4870 11090 4922
rect 14715 4870 14767 4922
rect 14779 4870 14831 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 12164 4768 12216 4820
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 15200 4768 15252 4820
rect 8668 4632 8720 4684
rect 12440 4700 12492 4752
rect 10140 4632 10192 4684
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 10416 4564 10468 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 11244 4564 11296 4616
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 11796 4564 11848 4616
rect 12164 4539 12216 4548
rect 8392 4428 8444 4480
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 12164 4505 12173 4539
rect 12173 4505 12207 4539
rect 12207 4505 12216 4539
rect 12164 4496 12216 4505
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14464 4564 14516 4616
rect 15108 4564 15160 4616
rect 13268 4496 13320 4548
rect 13820 4496 13872 4548
rect 12532 4428 12584 4480
rect 12624 4428 12676 4480
rect 16028 4428 16080 4480
rect 4882 4326 4934 4378
rect 4946 4326 4998 4378
rect 5010 4326 5062 4378
rect 5074 4326 5126 4378
rect 5138 4326 5190 4378
rect 8815 4326 8867 4378
rect 8879 4326 8931 4378
rect 8943 4326 8995 4378
rect 9007 4326 9059 4378
rect 9071 4326 9123 4378
rect 12748 4326 12800 4378
rect 12812 4326 12864 4378
rect 12876 4326 12928 4378
rect 12940 4326 12992 4378
rect 13004 4326 13056 4378
rect 16681 4326 16733 4378
rect 16745 4326 16797 4378
rect 16809 4326 16861 4378
rect 16873 4326 16925 4378
rect 16937 4326 16989 4378
rect 8484 4224 8536 4276
rect 12532 4224 12584 4276
rect 13176 4224 13228 4276
rect 13544 4224 13596 4276
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 8668 4088 8720 4140
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 9220 4020 9272 4072
rect 10140 4088 10192 4140
rect 11152 4088 11204 4140
rect 11796 4088 11848 4140
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 12808 4088 12860 4140
rect 13728 4088 13780 4140
rect 15292 4088 15344 4140
rect 15476 4088 15528 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 9680 4020 9732 4072
rect 10692 3952 10744 4004
rect 11612 3952 11664 4004
rect 8576 3884 8628 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 9680 3884 9732 3936
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12716 3884 12768 3936
rect 12808 3884 12860 3936
rect 13360 3884 13412 3936
rect 2916 3782 2968 3834
rect 2980 3782 3032 3834
rect 3044 3782 3096 3834
rect 3108 3782 3160 3834
rect 3172 3782 3224 3834
rect 6849 3782 6901 3834
rect 6913 3782 6965 3834
rect 6977 3782 7029 3834
rect 7041 3782 7093 3834
rect 7105 3782 7157 3834
rect 10782 3782 10834 3834
rect 10846 3782 10898 3834
rect 10910 3782 10962 3834
rect 10974 3782 11026 3834
rect 11038 3782 11090 3834
rect 14715 3782 14767 3834
rect 14779 3782 14831 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 11152 3680 11204 3732
rect 9312 3612 9364 3664
rect 11612 3680 11664 3732
rect 14280 3680 14332 3732
rect 13360 3612 13412 3664
rect 15108 3612 15160 3664
rect 11428 3544 11480 3596
rect 11980 3544 12032 3596
rect 12256 3476 12308 3528
rect 12624 3476 12676 3528
rect 12716 3476 12768 3528
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 16028 3519 16080 3528
rect 16028 3485 16046 3519
rect 16046 3485 16080 3519
rect 16028 3476 16080 3485
rect 16212 3476 16264 3528
rect 9220 3408 9272 3460
rect 11520 3408 11572 3460
rect 10416 3340 10468 3392
rect 11888 3383 11940 3392
rect 11888 3349 11897 3383
rect 11897 3349 11931 3383
rect 11931 3349 11940 3383
rect 11888 3340 11940 3349
rect 13176 3383 13228 3392
rect 13176 3349 13185 3383
rect 13185 3349 13219 3383
rect 13219 3349 13228 3383
rect 13176 3340 13228 3349
rect 16304 3340 16356 3392
rect 4882 3238 4934 3290
rect 4946 3238 4998 3290
rect 5010 3238 5062 3290
rect 5074 3238 5126 3290
rect 5138 3238 5190 3290
rect 8815 3238 8867 3290
rect 8879 3238 8931 3290
rect 8943 3238 8995 3290
rect 9007 3238 9059 3290
rect 9071 3238 9123 3290
rect 12748 3238 12800 3290
rect 12812 3238 12864 3290
rect 12876 3238 12928 3290
rect 12940 3238 12992 3290
rect 13004 3238 13056 3290
rect 16681 3238 16733 3290
rect 16745 3238 16797 3290
rect 16809 3238 16861 3290
rect 16873 3238 16925 3290
rect 16937 3238 16989 3290
rect 9220 3136 9272 3188
rect 13084 3136 13136 3188
rect 15476 3136 15528 3188
rect 11612 3068 11664 3120
rect 14556 3111 14608 3120
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 8208 3000 8260 3052
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 14556 3077 14565 3111
rect 14565 3077 14599 3111
rect 14599 3077 14608 3111
rect 14556 3068 14608 3077
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 13360 2864 13412 2916
rect 14464 2864 14516 2916
rect 8024 2839 8076 2848
rect 8024 2805 8033 2839
rect 8033 2805 8067 2839
rect 8067 2805 8076 2839
rect 8024 2796 8076 2805
rect 2916 2694 2968 2746
rect 2980 2694 3032 2746
rect 3044 2694 3096 2746
rect 3108 2694 3160 2746
rect 3172 2694 3224 2746
rect 6849 2694 6901 2746
rect 6913 2694 6965 2746
rect 6977 2694 7029 2746
rect 7041 2694 7093 2746
rect 7105 2694 7157 2746
rect 10782 2694 10834 2746
rect 10846 2694 10898 2746
rect 10910 2694 10962 2746
rect 10974 2694 11026 2746
rect 11038 2694 11090 2746
rect 14715 2694 14767 2746
rect 14779 2694 14831 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 8392 2592 8444 2644
rect 9404 2592 9456 2644
rect 10692 2592 10744 2644
rect 11704 2635 11756 2644
rect 11704 2601 11713 2635
rect 11713 2601 11747 2635
rect 11747 2601 11756 2635
rect 11704 2592 11756 2601
rect 12256 2592 12308 2644
rect 1584 2388 1636 2440
rect 4528 2388 4580 2440
rect 7472 2388 7524 2440
rect 8024 2388 8076 2440
rect 7748 2320 7800 2372
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 16212 2524 16264 2576
rect 8208 2388 8260 2397
rect 10416 2388 10468 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 13176 2388 13228 2440
rect 14556 2431 14608 2440
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 11428 2320 11480 2372
rect 12256 2252 12308 2304
rect 4882 2150 4934 2202
rect 4946 2150 4998 2202
rect 5010 2150 5062 2202
rect 5074 2150 5126 2202
rect 5138 2150 5190 2202
rect 8815 2150 8867 2202
rect 8879 2150 8931 2202
rect 8943 2150 8995 2202
rect 9007 2150 9059 2202
rect 9071 2150 9123 2202
rect 12748 2150 12800 2202
rect 12812 2150 12864 2202
rect 12876 2150 12928 2202
rect 12940 2150 12992 2202
rect 13004 2150 13056 2202
rect 16681 2150 16733 2202
rect 16745 2150 16797 2202
rect 16809 2150 16861 2202
rect 16873 2150 16925 2202
rect 16937 2150 16989 2202
<< metal2 >>
rect 1214 17200 1270 18000
rect 3422 17200 3478 18000
rect 5630 17354 5686 18000
rect 7838 17354 7894 18000
rect 10046 17354 10102 18000
rect 12254 17354 12310 18000
rect 5630 17326 5856 17354
rect 5630 17200 5686 17326
rect 1228 15706 1256 17200
rect 2916 15804 3224 15813
rect 2916 15802 2922 15804
rect 2978 15802 3002 15804
rect 3058 15802 3082 15804
rect 3138 15802 3162 15804
rect 3218 15802 3224 15804
rect 2978 15750 2980 15802
rect 3160 15750 3162 15802
rect 2916 15748 2922 15750
rect 2978 15748 3002 15750
rect 3058 15748 3082 15750
rect 3138 15748 3162 15750
rect 3218 15748 3224 15750
rect 2916 15739 3224 15748
rect 3436 15706 3464 17200
rect 5828 15706 5856 17326
rect 7838 17326 8064 17354
rect 7838 17200 7894 17326
rect 6849 15804 7157 15813
rect 6849 15802 6855 15804
rect 6911 15802 6935 15804
rect 6991 15802 7015 15804
rect 7071 15802 7095 15804
rect 7151 15802 7157 15804
rect 6911 15750 6913 15802
rect 7093 15750 7095 15802
rect 6849 15748 6855 15750
rect 6911 15748 6935 15750
rect 6991 15748 7015 15750
rect 7071 15748 7095 15750
rect 7151 15748 7157 15750
rect 6849 15739 7157 15748
rect 8036 15706 8064 17326
rect 10046 17326 10272 17354
rect 10046 17200 10102 17326
rect 10244 15706 10272 17326
rect 12254 17326 12388 17354
rect 12254 17200 12310 17326
rect 10782 15804 11090 15813
rect 10782 15802 10788 15804
rect 10844 15802 10868 15804
rect 10924 15802 10948 15804
rect 11004 15802 11028 15804
rect 11084 15802 11090 15804
rect 10844 15750 10846 15802
rect 11026 15750 11028 15802
rect 10782 15748 10788 15750
rect 10844 15748 10868 15750
rect 10924 15748 10948 15750
rect 11004 15748 11028 15750
rect 11084 15748 11090 15750
rect 10782 15739 11090 15748
rect 1216 15700 1268 15706
rect 1216 15642 1268 15648
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 10232 15700 10284 15706
rect 12360 15688 12388 17326
rect 14462 17200 14518 18000
rect 16670 17200 16726 18000
rect 14476 15706 14504 17200
rect 14715 15804 15023 15813
rect 14715 15802 14721 15804
rect 14777 15802 14801 15804
rect 14857 15802 14881 15804
rect 14937 15802 14961 15804
rect 15017 15802 15023 15804
rect 14777 15750 14779 15802
rect 14959 15750 14961 15802
rect 14715 15748 14721 15750
rect 14777 15748 14801 15750
rect 14857 15748 14881 15750
rect 14937 15748 14961 15750
rect 15017 15748 15023 15750
rect 14715 15739 15023 15748
rect 16684 15706 16712 17200
rect 12440 15700 12492 15706
rect 12360 15660 12440 15688
rect 10232 15642 10284 15648
rect 12440 15642 12492 15648
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 5574 2360 15302
rect 2916 14716 3224 14725
rect 2916 14714 2922 14716
rect 2978 14714 3002 14716
rect 3058 14714 3082 14716
rect 3138 14714 3162 14716
rect 3218 14714 3224 14716
rect 2978 14662 2980 14714
rect 3160 14662 3162 14714
rect 2916 14660 2922 14662
rect 2978 14660 3002 14662
rect 3058 14660 3082 14662
rect 3138 14660 3162 14662
rect 3218 14660 3224 14662
rect 2916 14651 3224 14660
rect 2916 13628 3224 13637
rect 2916 13626 2922 13628
rect 2978 13626 3002 13628
rect 3058 13626 3082 13628
rect 3138 13626 3162 13628
rect 3218 13626 3224 13628
rect 2978 13574 2980 13626
rect 3160 13574 3162 13626
rect 2916 13572 2922 13574
rect 2978 13572 3002 13574
rect 3058 13572 3082 13574
rect 3138 13572 3162 13574
rect 3218 13572 3224 13574
rect 2916 13563 3224 13572
rect 2916 12540 3224 12549
rect 2916 12538 2922 12540
rect 2978 12538 3002 12540
rect 3058 12538 3082 12540
rect 3138 12538 3162 12540
rect 3218 12538 3224 12540
rect 2978 12486 2980 12538
rect 3160 12486 3162 12538
rect 2916 12484 2922 12486
rect 2978 12484 3002 12486
rect 3058 12484 3082 12486
rect 3138 12484 3162 12486
rect 3218 12484 3224 12486
rect 2916 12475 3224 12484
rect 2916 11452 3224 11461
rect 2916 11450 2922 11452
rect 2978 11450 3002 11452
rect 3058 11450 3082 11452
rect 3138 11450 3162 11452
rect 3218 11450 3224 11452
rect 2978 11398 2980 11450
rect 3160 11398 3162 11450
rect 2916 11396 2922 11398
rect 2978 11396 3002 11398
rect 3058 11396 3082 11398
rect 3138 11396 3162 11398
rect 3218 11396 3224 11398
rect 2916 11387 3224 11396
rect 2916 10364 3224 10373
rect 2916 10362 2922 10364
rect 2978 10362 3002 10364
rect 3058 10362 3082 10364
rect 3138 10362 3162 10364
rect 3218 10362 3224 10364
rect 2978 10310 2980 10362
rect 3160 10310 3162 10362
rect 2916 10308 2922 10310
rect 2978 10308 3002 10310
rect 3058 10308 3082 10310
rect 3138 10308 3162 10310
rect 3218 10308 3224 10310
rect 2916 10299 3224 10308
rect 2916 9276 3224 9285
rect 2916 9274 2922 9276
rect 2978 9274 3002 9276
rect 3058 9274 3082 9276
rect 3138 9274 3162 9276
rect 3218 9274 3224 9276
rect 2978 9222 2980 9274
rect 3160 9222 3162 9274
rect 2916 9220 2922 9222
rect 2978 9220 3002 9222
rect 3058 9220 3082 9222
rect 3138 9220 3162 9222
rect 3218 9220 3224 9222
rect 2916 9211 3224 9220
rect 2916 8188 3224 8197
rect 2916 8186 2922 8188
rect 2978 8186 3002 8188
rect 3058 8186 3082 8188
rect 3138 8186 3162 8188
rect 3218 8186 3224 8188
rect 2978 8134 2980 8186
rect 3160 8134 3162 8186
rect 2916 8132 2922 8134
rect 2978 8132 3002 8134
rect 3058 8132 3082 8134
rect 3138 8132 3162 8134
rect 3218 8132 3224 8134
rect 2916 8123 3224 8132
rect 2916 7100 3224 7109
rect 2916 7098 2922 7100
rect 2978 7098 3002 7100
rect 3058 7098 3082 7100
rect 3138 7098 3162 7100
rect 3218 7098 3224 7100
rect 2978 7046 2980 7098
rect 3160 7046 3162 7098
rect 2916 7044 2922 7046
rect 2978 7044 3002 7046
rect 3058 7044 3082 7046
rect 3138 7044 3162 7046
rect 3218 7044 3224 7046
rect 2916 7035 3224 7044
rect 2916 6012 3224 6021
rect 2916 6010 2922 6012
rect 2978 6010 3002 6012
rect 3058 6010 3082 6012
rect 3138 6010 3162 6012
rect 3218 6010 3224 6012
rect 2978 5958 2980 6010
rect 3160 5958 3162 6010
rect 2916 5956 2922 5958
rect 2978 5956 3002 5958
rect 3058 5956 3082 5958
rect 3138 5956 3162 5958
rect 3218 5956 3224 5958
rect 2916 5947 3224 5956
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 4264 5370 4292 15438
rect 4882 15260 5190 15269
rect 4882 15258 4888 15260
rect 4944 15258 4968 15260
rect 5024 15258 5048 15260
rect 5104 15258 5128 15260
rect 5184 15258 5190 15260
rect 4944 15206 4946 15258
rect 5126 15206 5128 15258
rect 4882 15204 4888 15206
rect 4944 15204 4968 15206
rect 5024 15204 5048 15206
rect 5104 15204 5128 15206
rect 5184 15204 5190 15206
rect 4882 15195 5190 15204
rect 8815 15260 9123 15269
rect 8815 15258 8821 15260
rect 8877 15258 8901 15260
rect 8957 15258 8981 15260
rect 9037 15258 9061 15260
rect 9117 15258 9123 15260
rect 8877 15206 8879 15258
rect 9059 15206 9061 15258
rect 8815 15204 8821 15206
rect 8877 15204 8901 15206
rect 8957 15204 8981 15206
rect 9037 15204 9061 15206
rect 9117 15204 9123 15206
rect 8815 15195 9123 15204
rect 6849 14716 7157 14725
rect 6849 14714 6855 14716
rect 6911 14714 6935 14716
rect 6991 14714 7015 14716
rect 7071 14714 7095 14716
rect 7151 14714 7157 14716
rect 6911 14662 6913 14714
rect 7093 14662 7095 14714
rect 6849 14660 6855 14662
rect 6911 14660 6935 14662
rect 6991 14660 7015 14662
rect 7071 14660 7095 14662
rect 7151 14660 7157 14662
rect 6849 14651 7157 14660
rect 4882 14172 5190 14181
rect 4882 14170 4888 14172
rect 4944 14170 4968 14172
rect 5024 14170 5048 14172
rect 5104 14170 5128 14172
rect 5184 14170 5190 14172
rect 4944 14118 4946 14170
rect 5126 14118 5128 14170
rect 4882 14116 4888 14118
rect 4944 14116 4968 14118
rect 5024 14116 5048 14118
rect 5104 14116 5128 14118
rect 5184 14116 5190 14118
rect 4882 14107 5190 14116
rect 8815 14172 9123 14181
rect 8815 14170 8821 14172
rect 8877 14170 8901 14172
rect 8957 14170 8981 14172
rect 9037 14170 9061 14172
rect 9117 14170 9123 14172
rect 8877 14118 8879 14170
rect 9059 14118 9061 14170
rect 8815 14116 8821 14118
rect 8877 14116 8901 14118
rect 8957 14116 8981 14118
rect 9037 14116 9061 14118
rect 9117 14116 9123 14118
rect 8815 14107 9123 14116
rect 6849 13628 7157 13637
rect 6849 13626 6855 13628
rect 6911 13626 6935 13628
rect 6991 13626 7015 13628
rect 7071 13626 7095 13628
rect 7151 13626 7157 13628
rect 6911 13574 6913 13626
rect 7093 13574 7095 13626
rect 6849 13572 6855 13574
rect 6911 13572 6935 13574
rect 6991 13572 7015 13574
rect 7071 13572 7095 13574
rect 7151 13572 7157 13574
rect 6849 13563 7157 13572
rect 4882 13084 5190 13093
rect 4882 13082 4888 13084
rect 4944 13082 4968 13084
rect 5024 13082 5048 13084
rect 5104 13082 5128 13084
rect 5184 13082 5190 13084
rect 4944 13030 4946 13082
rect 5126 13030 5128 13082
rect 4882 13028 4888 13030
rect 4944 13028 4968 13030
rect 5024 13028 5048 13030
rect 5104 13028 5128 13030
rect 5184 13028 5190 13030
rect 4882 13019 5190 13028
rect 8815 13084 9123 13093
rect 8815 13082 8821 13084
rect 8877 13082 8901 13084
rect 8957 13082 8981 13084
rect 9037 13082 9061 13084
rect 9117 13082 9123 13084
rect 8877 13030 8879 13082
rect 9059 13030 9061 13082
rect 8815 13028 8821 13030
rect 8877 13028 8901 13030
rect 8957 13028 8981 13030
rect 9037 13028 9061 13030
rect 9117 13028 9123 13030
rect 8815 13019 9123 13028
rect 6849 12540 7157 12549
rect 6849 12538 6855 12540
rect 6911 12538 6935 12540
rect 6991 12538 7015 12540
rect 7071 12538 7095 12540
rect 7151 12538 7157 12540
rect 6911 12486 6913 12538
rect 7093 12486 7095 12538
rect 6849 12484 6855 12486
rect 6911 12484 6935 12486
rect 6991 12484 7015 12486
rect 7071 12484 7095 12486
rect 7151 12484 7157 12486
rect 6849 12475 7157 12484
rect 4882 11996 5190 12005
rect 4882 11994 4888 11996
rect 4944 11994 4968 11996
rect 5024 11994 5048 11996
rect 5104 11994 5128 11996
rect 5184 11994 5190 11996
rect 4944 11942 4946 11994
rect 5126 11942 5128 11994
rect 4882 11940 4888 11942
rect 4944 11940 4968 11942
rect 5024 11940 5048 11942
rect 5104 11940 5128 11942
rect 5184 11940 5190 11942
rect 4882 11931 5190 11940
rect 8815 11996 9123 12005
rect 8815 11994 8821 11996
rect 8877 11994 8901 11996
rect 8957 11994 8981 11996
rect 9037 11994 9061 11996
rect 9117 11994 9123 11996
rect 8877 11942 8879 11994
rect 9059 11942 9061 11994
rect 8815 11940 8821 11942
rect 8877 11940 8901 11942
rect 8957 11940 8981 11942
rect 9037 11940 9061 11942
rect 9117 11940 9123 11942
rect 8815 11931 9123 11940
rect 6849 11452 7157 11461
rect 6849 11450 6855 11452
rect 6911 11450 6935 11452
rect 6991 11450 7015 11452
rect 7071 11450 7095 11452
rect 7151 11450 7157 11452
rect 6911 11398 6913 11450
rect 7093 11398 7095 11450
rect 6849 11396 6855 11398
rect 6911 11396 6935 11398
rect 6991 11396 7015 11398
rect 7071 11396 7095 11398
rect 7151 11396 7157 11398
rect 6849 11387 7157 11396
rect 4882 10908 5190 10917
rect 4882 10906 4888 10908
rect 4944 10906 4968 10908
rect 5024 10906 5048 10908
rect 5104 10906 5128 10908
rect 5184 10906 5190 10908
rect 4944 10854 4946 10906
rect 5126 10854 5128 10906
rect 4882 10852 4888 10854
rect 4944 10852 4968 10854
rect 5024 10852 5048 10854
rect 5104 10852 5128 10854
rect 5184 10852 5190 10854
rect 4882 10843 5190 10852
rect 8815 10908 9123 10917
rect 8815 10906 8821 10908
rect 8877 10906 8901 10908
rect 8957 10906 8981 10908
rect 9037 10906 9061 10908
rect 9117 10906 9123 10908
rect 8877 10854 8879 10906
rect 9059 10854 9061 10906
rect 8815 10852 8821 10854
rect 8877 10852 8901 10854
rect 8957 10852 8981 10854
rect 9037 10852 9061 10854
rect 9117 10852 9123 10854
rect 8815 10843 9123 10852
rect 6849 10364 7157 10373
rect 6849 10362 6855 10364
rect 6911 10362 6935 10364
rect 6991 10362 7015 10364
rect 7071 10362 7095 10364
rect 7151 10362 7157 10364
rect 6911 10310 6913 10362
rect 7093 10310 7095 10362
rect 6849 10308 6855 10310
rect 6911 10308 6935 10310
rect 6991 10308 7015 10310
rect 7071 10308 7095 10310
rect 7151 10308 7157 10310
rect 6849 10299 7157 10308
rect 4882 9820 5190 9829
rect 4882 9818 4888 9820
rect 4944 9818 4968 9820
rect 5024 9818 5048 9820
rect 5104 9818 5128 9820
rect 5184 9818 5190 9820
rect 4944 9766 4946 9818
rect 5126 9766 5128 9818
rect 4882 9764 4888 9766
rect 4944 9764 4968 9766
rect 5024 9764 5048 9766
rect 5104 9764 5128 9766
rect 5184 9764 5190 9766
rect 4882 9755 5190 9764
rect 8815 9820 9123 9829
rect 8815 9818 8821 9820
rect 8877 9818 8901 9820
rect 8957 9818 8981 9820
rect 9037 9818 9061 9820
rect 9117 9818 9123 9820
rect 8877 9766 8879 9818
rect 9059 9766 9061 9818
rect 8815 9764 8821 9766
rect 8877 9764 8901 9766
rect 8957 9764 8981 9766
rect 9037 9764 9061 9766
rect 9117 9764 9123 9766
rect 8815 9755 9123 9764
rect 6849 9276 7157 9285
rect 6849 9274 6855 9276
rect 6911 9274 6935 9276
rect 6991 9274 7015 9276
rect 7071 9274 7095 9276
rect 7151 9274 7157 9276
rect 6911 9222 6913 9274
rect 7093 9222 7095 9274
rect 6849 9220 6855 9222
rect 6911 9220 6935 9222
rect 6991 9220 7015 9222
rect 7071 9220 7095 9222
rect 7151 9220 7157 9222
rect 6849 9211 7157 9220
rect 4882 8732 5190 8741
rect 4882 8730 4888 8732
rect 4944 8730 4968 8732
rect 5024 8730 5048 8732
rect 5104 8730 5128 8732
rect 5184 8730 5190 8732
rect 4944 8678 4946 8730
rect 5126 8678 5128 8730
rect 4882 8676 4888 8678
rect 4944 8676 4968 8678
rect 5024 8676 5048 8678
rect 5104 8676 5128 8678
rect 5184 8676 5190 8678
rect 4882 8667 5190 8676
rect 8815 8732 9123 8741
rect 8815 8730 8821 8732
rect 8877 8730 8901 8732
rect 8957 8730 8981 8732
rect 9037 8730 9061 8732
rect 9117 8730 9123 8732
rect 8877 8678 8879 8730
rect 9059 8678 9061 8730
rect 8815 8676 8821 8678
rect 8877 8676 8901 8678
rect 8957 8676 8981 8678
rect 9037 8676 9061 8678
rect 9117 8676 9123 8678
rect 8815 8667 9123 8676
rect 6849 8188 7157 8197
rect 6849 8186 6855 8188
rect 6911 8186 6935 8188
rect 6991 8186 7015 8188
rect 7071 8186 7095 8188
rect 7151 8186 7157 8188
rect 6911 8134 6913 8186
rect 7093 8134 7095 8186
rect 6849 8132 6855 8134
rect 6911 8132 6935 8134
rect 6991 8132 7015 8134
rect 7071 8132 7095 8134
rect 7151 8132 7157 8134
rect 6849 8123 7157 8132
rect 4882 7644 5190 7653
rect 4882 7642 4888 7644
rect 4944 7642 4968 7644
rect 5024 7642 5048 7644
rect 5104 7642 5128 7644
rect 5184 7642 5190 7644
rect 4944 7590 4946 7642
rect 5126 7590 5128 7642
rect 4882 7588 4888 7590
rect 4944 7588 4968 7590
rect 5024 7588 5048 7590
rect 5104 7588 5128 7590
rect 5184 7588 5190 7590
rect 4882 7579 5190 7588
rect 8815 7644 9123 7653
rect 8815 7642 8821 7644
rect 8877 7642 8901 7644
rect 8957 7642 8981 7644
rect 9037 7642 9061 7644
rect 9117 7642 9123 7644
rect 8877 7590 8879 7642
rect 9059 7590 9061 7642
rect 8815 7588 8821 7590
rect 8877 7588 8901 7590
rect 8957 7588 8981 7590
rect 9037 7588 9061 7590
rect 9117 7588 9123 7590
rect 8815 7579 9123 7588
rect 6849 7100 7157 7109
rect 6849 7098 6855 7100
rect 6911 7098 6935 7100
rect 6991 7098 7015 7100
rect 7071 7098 7095 7100
rect 7151 7098 7157 7100
rect 6911 7046 6913 7098
rect 7093 7046 7095 7098
rect 6849 7044 6855 7046
rect 6911 7044 6935 7046
rect 6991 7044 7015 7046
rect 7071 7044 7095 7046
rect 7151 7044 7157 7046
rect 6849 7035 7157 7044
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 4882 6556 5190 6565
rect 4882 6554 4888 6556
rect 4944 6554 4968 6556
rect 5024 6554 5048 6556
rect 5104 6554 5128 6556
rect 5184 6554 5190 6556
rect 4944 6502 4946 6554
rect 5126 6502 5128 6554
rect 4882 6500 4888 6502
rect 4944 6500 4968 6502
rect 5024 6500 5048 6502
rect 5104 6500 5128 6502
rect 5184 6500 5190 6502
rect 4882 6491 5190 6500
rect 8815 6556 9123 6565
rect 8815 6554 8821 6556
rect 8877 6554 8901 6556
rect 8957 6554 8981 6556
rect 9037 6554 9061 6556
rect 9117 6554 9123 6556
rect 8877 6502 8879 6554
rect 9059 6502 9061 6554
rect 8815 6500 8821 6502
rect 8877 6500 8901 6502
rect 8957 6500 8981 6502
rect 9037 6500 9061 6502
rect 9117 6500 9123 6502
rect 8815 6491 9123 6500
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 6849 6012 7157 6021
rect 6849 6010 6855 6012
rect 6911 6010 6935 6012
rect 6991 6010 7015 6012
rect 7071 6010 7095 6012
rect 7151 6010 7157 6012
rect 6911 5958 6913 6010
rect 7093 5958 7095 6010
rect 6849 5956 6855 5958
rect 6911 5956 6935 5958
rect 6991 5956 7015 5958
rect 7071 5956 7095 5958
rect 7151 5956 7157 5958
rect 6849 5947 7157 5956
rect 9140 5778 9168 6054
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 4882 5468 5190 5477
rect 4882 5466 4888 5468
rect 4944 5466 4968 5468
rect 5024 5466 5048 5468
rect 5104 5466 5128 5468
rect 5184 5466 5190 5468
rect 4944 5414 4946 5466
rect 5126 5414 5128 5466
rect 4882 5412 4888 5414
rect 4944 5412 4968 5414
rect 5024 5412 5048 5414
rect 5104 5412 5128 5414
rect 5184 5412 5190 5414
rect 4882 5403 5190 5412
rect 8815 5468 9123 5477
rect 8815 5466 8821 5468
rect 8877 5466 8901 5468
rect 8957 5466 8981 5468
rect 9037 5466 9061 5468
rect 9117 5466 9123 5468
rect 8877 5414 8879 5466
rect 9059 5414 9061 5466
rect 8815 5412 8821 5414
rect 8877 5412 8901 5414
rect 8957 5412 8981 5414
rect 9037 5412 9061 5414
rect 9117 5412 9123 5414
rect 8815 5403 9123 5412
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 2916 4924 3224 4933
rect 2916 4922 2922 4924
rect 2978 4922 3002 4924
rect 3058 4922 3082 4924
rect 3138 4922 3162 4924
rect 3218 4922 3224 4924
rect 2978 4870 2980 4922
rect 3160 4870 3162 4922
rect 2916 4868 2922 4870
rect 2978 4868 3002 4870
rect 3058 4868 3082 4870
rect 3138 4868 3162 4870
rect 3218 4868 3224 4870
rect 2916 4859 3224 4868
rect 6849 4924 7157 4933
rect 6849 4922 6855 4924
rect 6911 4922 6935 4924
rect 6991 4922 7015 4924
rect 7071 4922 7095 4924
rect 7151 4922 7157 4924
rect 6911 4870 6913 4922
rect 7093 4870 7095 4922
rect 6849 4868 6855 4870
rect 6911 4868 6935 4870
rect 6991 4868 7015 4870
rect 7071 4868 7095 4870
rect 7151 4868 7157 4870
rect 6849 4859 7157 4868
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 4882 4380 5190 4389
rect 4882 4378 4888 4380
rect 4944 4378 4968 4380
rect 5024 4378 5048 4380
rect 5104 4378 5128 4380
rect 5184 4378 5190 4380
rect 4944 4326 4946 4378
rect 5126 4326 5128 4378
rect 4882 4324 4888 4326
rect 4944 4324 4968 4326
rect 5024 4324 5048 4326
rect 5104 4324 5128 4326
rect 5184 4324 5190 4326
rect 4882 4315 5190 4324
rect 8404 4146 8432 4422
rect 8496 4282 8524 5102
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8588 3942 8616 4762
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4146 8708 4626
rect 8815 4380 9123 4389
rect 8815 4378 8821 4380
rect 8877 4378 8901 4380
rect 8957 4378 8981 4380
rect 9037 4378 9061 4380
rect 9117 4378 9123 4380
rect 8877 4326 8879 4378
rect 9059 4326 9061 4378
rect 8815 4324 8821 4326
rect 8877 4324 8901 4326
rect 8957 4324 8981 4326
rect 9037 4324 9061 4326
rect 9117 4324 9123 4326
rect 8815 4315 9123 4324
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 9232 4078 9260 6258
rect 9416 5710 9444 6326
rect 9876 6322 9904 6598
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 10152 5914 10180 15438
rect 10704 6118 10732 15506
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 12748 15260 13056 15269
rect 12748 15258 12754 15260
rect 12810 15258 12834 15260
rect 12890 15258 12914 15260
rect 12970 15258 12994 15260
rect 13050 15258 13056 15260
rect 12810 15206 12812 15258
rect 12992 15206 12994 15258
rect 12748 15204 12754 15206
rect 12810 15204 12834 15206
rect 12890 15204 12914 15206
rect 12970 15204 12994 15206
rect 13050 15204 13056 15206
rect 12748 15195 13056 15204
rect 10782 14716 11090 14725
rect 10782 14714 10788 14716
rect 10844 14714 10868 14716
rect 10924 14714 10948 14716
rect 11004 14714 11028 14716
rect 11084 14714 11090 14716
rect 10844 14662 10846 14714
rect 11026 14662 11028 14714
rect 10782 14660 10788 14662
rect 10844 14660 10868 14662
rect 10924 14660 10948 14662
rect 11004 14660 11028 14662
rect 11084 14660 11090 14662
rect 10782 14651 11090 14660
rect 12748 14172 13056 14181
rect 12748 14170 12754 14172
rect 12810 14170 12834 14172
rect 12890 14170 12914 14172
rect 12970 14170 12994 14172
rect 13050 14170 13056 14172
rect 12810 14118 12812 14170
rect 12992 14118 12994 14170
rect 12748 14116 12754 14118
rect 12810 14116 12834 14118
rect 12890 14116 12914 14118
rect 12970 14116 12994 14118
rect 13050 14116 13056 14118
rect 12748 14107 13056 14116
rect 10782 13628 11090 13637
rect 10782 13626 10788 13628
rect 10844 13626 10868 13628
rect 10924 13626 10948 13628
rect 11004 13626 11028 13628
rect 11084 13626 11090 13628
rect 10844 13574 10846 13626
rect 11026 13574 11028 13626
rect 10782 13572 10788 13574
rect 10844 13572 10868 13574
rect 10924 13572 10948 13574
rect 11004 13572 11028 13574
rect 11084 13572 11090 13574
rect 10782 13563 11090 13572
rect 12748 13084 13056 13093
rect 12748 13082 12754 13084
rect 12810 13082 12834 13084
rect 12890 13082 12914 13084
rect 12970 13082 12994 13084
rect 13050 13082 13056 13084
rect 12810 13030 12812 13082
rect 12992 13030 12994 13082
rect 12748 13028 12754 13030
rect 12810 13028 12834 13030
rect 12890 13028 12914 13030
rect 12970 13028 12994 13030
rect 13050 13028 13056 13030
rect 12748 13019 13056 13028
rect 10782 12540 11090 12549
rect 10782 12538 10788 12540
rect 10844 12538 10868 12540
rect 10924 12538 10948 12540
rect 11004 12538 11028 12540
rect 11084 12538 11090 12540
rect 10844 12486 10846 12538
rect 11026 12486 11028 12538
rect 10782 12484 10788 12486
rect 10844 12484 10868 12486
rect 10924 12484 10948 12486
rect 11004 12484 11028 12486
rect 11084 12484 11090 12486
rect 10782 12475 11090 12484
rect 12748 11996 13056 12005
rect 12748 11994 12754 11996
rect 12810 11994 12834 11996
rect 12890 11994 12914 11996
rect 12970 11994 12994 11996
rect 13050 11994 13056 11996
rect 12810 11942 12812 11994
rect 12992 11942 12994 11994
rect 12748 11940 12754 11942
rect 12810 11940 12834 11942
rect 12890 11940 12914 11942
rect 12970 11940 12994 11942
rect 13050 11940 13056 11942
rect 12748 11931 13056 11940
rect 10782 11452 11090 11461
rect 10782 11450 10788 11452
rect 10844 11450 10868 11452
rect 10924 11450 10948 11452
rect 11004 11450 11028 11452
rect 11084 11450 11090 11452
rect 10844 11398 10846 11450
rect 11026 11398 11028 11450
rect 10782 11396 10788 11398
rect 10844 11396 10868 11398
rect 10924 11396 10948 11398
rect 11004 11396 11028 11398
rect 11084 11396 11090 11398
rect 10782 11387 11090 11396
rect 12748 10908 13056 10917
rect 12748 10906 12754 10908
rect 12810 10906 12834 10908
rect 12890 10906 12914 10908
rect 12970 10906 12994 10908
rect 13050 10906 13056 10908
rect 12810 10854 12812 10906
rect 12992 10854 12994 10906
rect 12748 10852 12754 10854
rect 12810 10852 12834 10854
rect 12890 10852 12914 10854
rect 12970 10852 12994 10854
rect 13050 10852 13056 10854
rect 12748 10843 13056 10852
rect 10782 10364 11090 10373
rect 10782 10362 10788 10364
rect 10844 10362 10868 10364
rect 10924 10362 10948 10364
rect 11004 10362 11028 10364
rect 11084 10362 11090 10364
rect 10844 10310 10846 10362
rect 11026 10310 11028 10362
rect 10782 10308 10788 10310
rect 10844 10308 10868 10310
rect 10924 10308 10948 10310
rect 11004 10308 11028 10310
rect 11084 10308 11090 10310
rect 10782 10299 11090 10308
rect 12748 9820 13056 9829
rect 12748 9818 12754 9820
rect 12810 9818 12834 9820
rect 12890 9818 12914 9820
rect 12970 9818 12994 9820
rect 13050 9818 13056 9820
rect 12810 9766 12812 9818
rect 12992 9766 12994 9818
rect 12748 9764 12754 9766
rect 12810 9764 12834 9766
rect 12890 9764 12914 9766
rect 12970 9764 12994 9766
rect 13050 9764 13056 9766
rect 12748 9755 13056 9764
rect 10782 9276 11090 9285
rect 10782 9274 10788 9276
rect 10844 9274 10868 9276
rect 10924 9274 10948 9276
rect 11004 9274 11028 9276
rect 11084 9274 11090 9276
rect 10844 9222 10846 9274
rect 11026 9222 11028 9274
rect 10782 9220 10788 9222
rect 10844 9220 10868 9222
rect 10924 9220 10948 9222
rect 11004 9220 11028 9222
rect 11084 9220 11090 9222
rect 10782 9211 11090 9220
rect 12748 8732 13056 8741
rect 12748 8730 12754 8732
rect 12810 8730 12834 8732
rect 12890 8730 12914 8732
rect 12970 8730 12994 8732
rect 13050 8730 13056 8732
rect 12810 8678 12812 8730
rect 12992 8678 12994 8730
rect 12748 8676 12754 8678
rect 12810 8676 12834 8678
rect 12890 8676 12914 8678
rect 12970 8676 12994 8678
rect 13050 8676 13056 8678
rect 12748 8667 13056 8676
rect 10782 8188 11090 8197
rect 10782 8186 10788 8188
rect 10844 8186 10868 8188
rect 10924 8186 10948 8188
rect 11004 8186 11028 8188
rect 11084 8186 11090 8188
rect 10844 8134 10846 8186
rect 11026 8134 11028 8186
rect 10782 8132 10788 8134
rect 10844 8132 10868 8134
rect 10924 8132 10948 8134
rect 11004 8132 11028 8134
rect 11084 8132 11090 8134
rect 10782 8123 11090 8132
rect 12748 7644 13056 7653
rect 12748 7642 12754 7644
rect 12810 7642 12834 7644
rect 12890 7642 12914 7644
rect 12970 7642 12994 7644
rect 13050 7642 13056 7644
rect 12810 7590 12812 7642
rect 12992 7590 12994 7642
rect 12748 7588 12754 7590
rect 12810 7588 12834 7590
rect 12890 7588 12914 7590
rect 12970 7588 12994 7590
rect 13050 7588 13056 7590
rect 12748 7579 13056 7588
rect 10782 7100 11090 7109
rect 10782 7098 10788 7100
rect 10844 7098 10868 7100
rect 10924 7098 10948 7100
rect 11004 7098 11028 7100
rect 11084 7098 11090 7100
rect 10844 7046 10846 7098
rect 11026 7046 11028 7098
rect 10782 7044 10788 7046
rect 10844 7044 10868 7046
rect 10924 7044 10948 7046
rect 11004 7044 11028 7046
rect 11084 7044 11090 7046
rect 10782 7035 11090 7044
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 5234 9444 5646
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9508 4622 9536 5306
rect 10152 4690 10180 5850
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10428 4622 10456 6054
rect 10782 6012 11090 6021
rect 10782 6010 10788 6012
rect 10844 6010 10868 6012
rect 10924 6010 10948 6012
rect 11004 6010 11028 6012
rect 11084 6010 11090 6012
rect 10844 5958 10846 6010
rect 11026 5958 11028 6010
rect 10782 5956 10788 5958
rect 10844 5956 10868 5958
rect 10924 5956 10948 5958
rect 11004 5956 11028 5958
rect 11084 5956 11090 5958
rect 10782 5947 11090 5956
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11256 5658 11284 6734
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 5914 11376 6190
rect 12636 5914 12664 6734
rect 12748 6556 13056 6565
rect 12748 6554 12754 6556
rect 12810 6554 12834 6556
rect 12890 6554 12914 6556
rect 12970 6554 12994 6556
rect 13050 6554 13056 6556
rect 12810 6502 12812 6554
rect 12992 6502 12994 6554
rect 12748 6500 12754 6502
rect 12810 6500 12834 6502
rect 12890 6500 12914 6502
rect 12970 6500 12994 6502
rect 13050 6500 13056 6502
rect 12748 6491 13056 6500
rect 13188 6118 13216 15438
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13648 6662 13676 15370
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13280 5914 13308 6190
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 11164 5370 11192 5646
rect 11256 5630 11376 5658
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10782 4924 11090 4933
rect 10782 4922 10788 4924
rect 10844 4922 10868 4924
rect 10924 4922 10948 4924
rect 11004 4922 11028 4924
rect 11084 4922 11090 4924
rect 10844 4870 10846 4922
rect 11026 4870 11028 4922
rect 10782 4868 10788 4870
rect 10844 4868 10868 4870
rect 10924 4868 10948 4870
rect 11004 4868 11028 4870
rect 11084 4868 11090 4870
rect 10782 4859 11090 4868
rect 11256 4622 11284 5510
rect 11348 4826 11376 5630
rect 12360 5098 12388 5714
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 2916 3836 3224 3845
rect 2916 3834 2922 3836
rect 2978 3834 3002 3836
rect 3058 3834 3082 3836
rect 3138 3834 3162 3836
rect 3218 3834 3224 3836
rect 2978 3782 2980 3834
rect 3160 3782 3162 3834
rect 2916 3780 2922 3782
rect 2978 3780 3002 3782
rect 3058 3780 3082 3782
rect 3138 3780 3162 3782
rect 3218 3780 3224 3782
rect 2916 3771 3224 3780
rect 6849 3836 7157 3845
rect 6849 3834 6855 3836
rect 6911 3834 6935 3836
rect 6991 3834 7015 3836
rect 7071 3834 7095 3836
rect 7151 3834 7157 3836
rect 6911 3782 6913 3834
rect 7093 3782 7095 3834
rect 6849 3780 6855 3782
rect 6911 3780 6935 3782
rect 6991 3780 7015 3782
rect 7071 3780 7095 3782
rect 7151 3780 7157 3782
rect 6849 3771 7157 3780
rect 9232 3466 9260 3878
rect 9324 3670 9352 4082
rect 9692 4078 9720 4422
rect 10152 4146 10180 4422
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 10704 4010 10732 4558
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 4882 3292 5190 3301
rect 4882 3290 4888 3292
rect 4944 3290 4968 3292
rect 5024 3290 5048 3292
rect 5104 3290 5128 3292
rect 5184 3290 5190 3292
rect 4944 3238 4946 3290
rect 5126 3238 5128 3290
rect 4882 3236 4888 3238
rect 4944 3236 4968 3238
rect 5024 3236 5048 3238
rect 5104 3236 5128 3238
rect 5184 3236 5190 3238
rect 4882 3227 5190 3236
rect 8815 3292 9123 3301
rect 8815 3290 8821 3292
rect 8877 3290 8901 3292
rect 8957 3290 8981 3292
rect 9037 3290 9061 3292
rect 9117 3290 9123 3292
rect 8877 3238 8879 3290
rect 9059 3238 9061 3290
rect 8815 3236 8821 3238
rect 8877 3236 8901 3238
rect 8957 3236 8981 3238
rect 9037 3236 9061 3238
rect 9117 3236 9123 3238
rect 8815 3227 9123 3236
rect 9232 3194 9260 3402
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9692 3058 9720 3878
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 2916 2748 3224 2757
rect 2916 2746 2922 2748
rect 2978 2746 3002 2748
rect 3058 2746 3082 2748
rect 3138 2746 3162 2748
rect 3218 2746 3224 2748
rect 2978 2694 2980 2746
rect 3160 2694 3162 2746
rect 2916 2692 2922 2694
rect 2978 2692 3002 2694
rect 3058 2692 3082 2694
rect 3138 2692 3162 2694
rect 3218 2692 3224 2694
rect 2916 2683 3224 2692
rect 6849 2748 7157 2757
rect 6849 2746 6855 2748
rect 6911 2746 6935 2748
rect 6991 2746 7015 2748
rect 7071 2746 7095 2748
rect 7151 2746 7157 2748
rect 6911 2694 6913 2746
rect 7093 2694 7095 2746
rect 6849 2692 6855 2694
rect 6911 2692 6935 2694
rect 6991 2692 7015 2694
rect 7071 2692 7095 2694
rect 7151 2692 7157 2694
rect 6849 2683 7157 2692
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 1596 800 1624 2382
rect 4540 800 4568 2382
rect 4882 2204 5190 2213
rect 4882 2202 4888 2204
rect 4944 2202 4968 2204
rect 5024 2202 5048 2204
rect 5104 2202 5128 2204
rect 5184 2202 5190 2204
rect 4944 2150 4946 2202
rect 5126 2150 5128 2202
rect 4882 2148 4888 2150
rect 4944 2148 4968 2150
rect 5024 2148 5048 2150
rect 5104 2148 5128 2150
rect 5184 2148 5190 2150
rect 4882 2139 5190 2148
rect 7484 800 7512 2382
rect 7760 2378 7788 2994
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8036 2446 8064 2790
rect 8220 2446 8248 2994
rect 8404 2650 8432 2994
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9416 2650 9444 2926
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 10428 2446 10456 3334
rect 10704 2650 10732 3946
rect 10782 3836 11090 3845
rect 10782 3834 10788 3836
rect 10844 3834 10868 3836
rect 10924 3834 10948 3836
rect 11004 3834 11028 3836
rect 11084 3834 11090 3836
rect 10844 3782 10846 3834
rect 11026 3782 11028 3834
rect 10782 3780 10788 3782
rect 10844 3780 10868 3782
rect 10924 3780 10948 3782
rect 11004 3780 11028 3782
rect 11084 3780 11090 3782
rect 10782 3771 11090 3780
rect 11164 3738 11192 4082
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 10782 2748 11090 2757
rect 10782 2746 10788 2748
rect 10844 2746 10868 2748
rect 10924 2746 10948 2748
rect 11004 2746 11028 2748
rect 11084 2746 11090 2748
rect 10844 2694 10846 2746
rect 11026 2694 11028 2746
rect 10782 2692 10788 2694
rect 10844 2692 10868 2694
rect 10924 2692 10948 2694
rect 11004 2692 11028 2694
rect 11084 2692 11090 2694
rect 10782 2683 11090 2692
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 8815 2204 9123 2213
rect 8815 2202 8821 2204
rect 8877 2202 8901 2204
rect 8957 2202 8981 2204
rect 9037 2202 9061 2204
rect 9117 2202 9123 2204
rect 8877 2150 8879 2202
rect 9059 2150 9061 2202
rect 8815 2148 8821 2150
rect 8877 2148 8901 2150
rect 8957 2148 8981 2150
rect 9037 2148 9061 2150
rect 9117 2148 9123 2150
rect 8815 2139 9123 2148
rect 10428 800 10456 2382
rect 11440 2378 11468 3538
rect 11532 3466 11560 4762
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11624 4010 11652 4558
rect 11808 4146 11836 4558
rect 12176 4554 12204 4762
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12360 4162 12388 5034
rect 12452 4758 12480 5102
rect 12544 4826 12572 5170
rect 12636 5030 12664 5714
rect 13556 5710 13584 6054
rect 13648 5778 13676 6598
rect 13740 6322 13768 6734
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13740 6202 13768 6258
rect 13740 6174 13860 6202
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 12748 5468 13056 5477
rect 12748 5466 12754 5468
rect 12810 5466 12834 5468
rect 12890 5466 12914 5468
rect 12970 5466 12994 5468
rect 13050 5466 13056 5468
rect 12810 5414 12812 5466
rect 12992 5414 12994 5466
rect 12748 5412 12754 5414
rect 12810 5412 12834 5414
rect 12890 5412 12914 5414
rect 12970 5412 12994 5414
rect 13050 5412 13056 5414
rect 12748 5403 13056 5412
rect 13096 5370 13124 5646
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12268 4134 12388 4162
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11624 3738 11652 3946
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11624 3126 11652 3674
rect 11992 3602 12020 4082
rect 12268 3942 12296 4134
rect 12452 3942 12480 4694
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12624 4480 12676 4486
rect 13188 4434 13216 5578
rect 13464 5370 13492 5646
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13268 4548 13320 4554
rect 13268 4490 13320 4496
rect 12624 4422 12676 4428
rect 12544 4282 12572 4422
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 12268 3534 12296 3878
rect 12636 3534 12664 4422
rect 13096 4406 13216 4434
rect 12748 4380 13056 4389
rect 12748 4378 12754 4380
rect 12810 4378 12834 4380
rect 12890 4378 12914 4380
rect 12970 4378 12994 4380
rect 13050 4378 13056 4380
rect 12810 4326 12812 4378
rect 12992 4326 12994 4378
rect 12748 4324 12754 4326
rect 12810 4324 12834 4326
rect 12890 4324 12914 4326
rect 12970 4324 12994 4326
rect 13050 4324 13056 4326
rect 12748 4315 13056 4324
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12820 3942 12848 4082
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12728 3534 12756 3878
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11716 2650 11744 2926
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11900 2446 11928 3334
rect 12268 2650 12296 3470
rect 12748 3292 13056 3301
rect 12748 3290 12754 3292
rect 12810 3290 12834 3292
rect 12890 3290 12914 3292
rect 12970 3290 12994 3292
rect 13050 3290 13056 3292
rect 12810 3238 12812 3290
rect 12992 3238 12994 3290
rect 12748 3236 12754 3238
rect 12810 3236 12834 3238
rect 12890 3236 12914 3238
rect 12970 3236 12994 3238
rect 13050 3236 13056 3238
rect 12748 3227 13056 3236
rect 13096 3194 13124 4406
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13188 3534 13216 4218
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11428 2372 11480 2378
rect 11428 2314 11480 2320
rect 12268 2310 12296 2586
rect 13188 2446 13216 3334
rect 13280 2990 13308 4490
rect 13372 3942 13400 4966
rect 13556 4282 13584 5170
rect 13740 5166 13768 5850
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13740 4146 13768 5102
rect 13832 4554 13860 6174
rect 14292 6118 14320 15438
rect 14715 14716 15023 14725
rect 14715 14714 14721 14716
rect 14777 14714 14801 14716
rect 14857 14714 14881 14716
rect 14937 14714 14961 14716
rect 15017 14714 15023 14716
rect 14777 14662 14779 14714
rect 14959 14662 14961 14714
rect 14715 14660 14721 14662
rect 14777 14660 14801 14662
rect 14857 14660 14881 14662
rect 14937 14660 14961 14662
rect 15017 14660 15023 14662
rect 14715 14651 15023 14660
rect 14715 13628 15023 13637
rect 14715 13626 14721 13628
rect 14777 13626 14801 13628
rect 14857 13626 14881 13628
rect 14937 13626 14961 13628
rect 15017 13626 15023 13628
rect 14777 13574 14779 13626
rect 14959 13574 14961 13626
rect 14715 13572 14721 13574
rect 14777 13572 14801 13574
rect 14857 13572 14881 13574
rect 14937 13572 14961 13574
rect 15017 13572 15023 13574
rect 14715 13563 15023 13572
rect 14715 12540 15023 12549
rect 14715 12538 14721 12540
rect 14777 12538 14801 12540
rect 14857 12538 14881 12540
rect 14937 12538 14961 12540
rect 15017 12538 15023 12540
rect 14777 12486 14779 12538
rect 14959 12486 14961 12538
rect 14715 12484 14721 12486
rect 14777 12484 14801 12486
rect 14857 12484 14881 12486
rect 14937 12484 14961 12486
rect 15017 12484 15023 12486
rect 14715 12475 15023 12484
rect 14715 11452 15023 11461
rect 14715 11450 14721 11452
rect 14777 11450 14801 11452
rect 14857 11450 14881 11452
rect 14937 11450 14961 11452
rect 15017 11450 15023 11452
rect 14777 11398 14779 11450
rect 14959 11398 14961 11450
rect 14715 11396 14721 11398
rect 14777 11396 14801 11398
rect 14857 11396 14881 11398
rect 14937 11396 14961 11398
rect 15017 11396 15023 11398
rect 14715 11387 15023 11396
rect 14715 10364 15023 10373
rect 14715 10362 14721 10364
rect 14777 10362 14801 10364
rect 14857 10362 14881 10364
rect 14937 10362 14961 10364
rect 15017 10362 15023 10364
rect 14777 10310 14779 10362
rect 14959 10310 14961 10362
rect 14715 10308 14721 10310
rect 14777 10308 14801 10310
rect 14857 10308 14881 10310
rect 14937 10308 14961 10310
rect 15017 10308 15023 10310
rect 14715 10299 15023 10308
rect 14715 9276 15023 9285
rect 14715 9274 14721 9276
rect 14777 9274 14801 9276
rect 14857 9274 14881 9276
rect 14937 9274 14961 9276
rect 15017 9274 15023 9276
rect 14777 9222 14779 9274
rect 14959 9222 14961 9274
rect 14715 9220 14721 9222
rect 14777 9220 14801 9222
rect 14857 9220 14881 9222
rect 14937 9220 14961 9222
rect 15017 9220 15023 9222
rect 14715 9211 15023 9220
rect 14715 8188 15023 8197
rect 14715 8186 14721 8188
rect 14777 8186 14801 8188
rect 14857 8186 14881 8188
rect 14937 8186 14961 8188
rect 15017 8186 15023 8188
rect 14777 8134 14779 8186
rect 14959 8134 14961 8186
rect 14715 8132 14721 8134
rect 14777 8132 14801 8134
rect 14857 8132 14881 8134
rect 14937 8132 14961 8134
rect 15017 8132 15023 8134
rect 14715 8123 15023 8132
rect 14715 7100 15023 7109
rect 14715 7098 14721 7100
rect 14777 7098 14801 7100
rect 14857 7098 14881 7100
rect 14937 7098 14961 7100
rect 15017 7098 15023 7100
rect 14777 7046 14779 7098
rect 14959 7046 14961 7098
rect 14715 7044 14721 7046
rect 14777 7044 14801 7046
rect 14857 7044 14881 7046
rect 14937 7044 14961 7046
rect 15017 7044 15023 7046
rect 14715 7035 15023 7044
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14715 6012 15023 6021
rect 14715 6010 14721 6012
rect 14777 6010 14801 6012
rect 14857 6010 14881 6012
rect 14937 6010 14961 6012
rect 15017 6010 15023 6012
rect 14777 5958 14779 6010
rect 14959 5958 14961 6010
rect 14715 5956 14721 5958
rect 14777 5956 14801 5958
rect 14857 5956 14881 5958
rect 14937 5956 14961 5958
rect 15017 5956 15023 5958
rect 14715 5947 15023 5956
rect 15212 5778 15240 15438
rect 16681 15260 16989 15269
rect 16681 15258 16687 15260
rect 16743 15258 16767 15260
rect 16823 15258 16847 15260
rect 16903 15258 16927 15260
rect 16983 15258 16989 15260
rect 16743 15206 16745 15258
rect 16925 15206 16927 15258
rect 16681 15204 16687 15206
rect 16743 15204 16767 15206
rect 16823 15204 16847 15206
rect 16903 15204 16927 15206
rect 16983 15204 16989 15206
rect 16681 15195 16989 15204
rect 16681 14172 16989 14181
rect 16681 14170 16687 14172
rect 16743 14170 16767 14172
rect 16823 14170 16847 14172
rect 16903 14170 16927 14172
rect 16983 14170 16989 14172
rect 16743 14118 16745 14170
rect 16925 14118 16927 14170
rect 16681 14116 16687 14118
rect 16743 14116 16767 14118
rect 16823 14116 16847 14118
rect 16903 14116 16927 14118
rect 16983 14116 16989 14118
rect 16681 14107 16989 14116
rect 16681 13084 16989 13093
rect 16681 13082 16687 13084
rect 16743 13082 16767 13084
rect 16823 13082 16847 13084
rect 16903 13082 16927 13084
rect 16983 13082 16989 13084
rect 16743 13030 16745 13082
rect 16925 13030 16927 13082
rect 16681 13028 16687 13030
rect 16743 13028 16767 13030
rect 16823 13028 16847 13030
rect 16903 13028 16927 13030
rect 16983 13028 16989 13030
rect 16681 13019 16989 13028
rect 16681 11996 16989 12005
rect 16681 11994 16687 11996
rect 16743 11994 16767 11996
rect 16823 11994 16847 11996
rect 16903 11994 16927 11996
rect 16983 11994 16989 11996
rect 16743 11942 16745 11994
rect 16925 11942 16927 11994
rect 16681 11940 16687 11942
rect 16743 11940 16767 11942
rect 16823 11940 16847 11942
rect 16903 11940 16927 11942
rect 16983 11940 16989 11942
rect 16681 11931 16989 11940
rect 16681 10908 16989 10917
rect 16681 10906 16687 10908
rect 16743 10906 16767 10908
rect 16823 10906 16847 10908
rect 16903 10906 16927 10908
rect 16983 10906 16989 10908
rect 16743 10854 16745 10906
rect 16925 10854 16927 10906
rect 16681 10852 16687 10854
rect 16743 10852 16767 10854
rect 16823 10852 16847 10854
rect 16903 10852 16927 10854
rect 16983 10852 16989 10854
rect 16681 10843 16989 10852
rect 16681 9820 16989 9829
rect 16681 9818 16687 9820
rect 16743 9818 16767 9820
rect 16823 9818 16847 9820
rect 16903 9818 16927 9820
rect 16983 9818 16989 9820
rect 16743 9766 16745 9818
rect 16925 9766 16927 9818
rect 16681 9764 16687 9766
rect 16743 9764 16767 9766
rect 16823 9764 16847 9766
rect 16903 9764 16927 9766
rect 16983 9764 16989 9766
rect 16681 9755 16989 9764
rect 16681 8732 16989 8741
rect 16681 8730 16687 8732
rect 16743 8730 16767 8732
rect 16823 8730 16847 8732
rect 16903 8730 16927 8732
rect 16983 8730 16989 8732
rect 16743 8678 16745 8730
rect 16925 8678 16927 8730
rect 16681 8676 16687 8678
rect 16743 8676 16767 8678
rect 16823 8676 16847 8678
rect 16903 8676 16927 8678
rect 16983 8676 16989 8678
rect 16681 8667 16989 8676
rect 16681 7644 16989 7653
rect 16681 7642 16687 7644
rect 16743 7642 16767 7644
rect 16823 7642 16847 7644
rect 16903 7642 16927 7644
rect 16983 7642 16989 7644
rect 16743 7590 16745 7642
rect 16925 7590 16927 7642
rect 16681 7588 16687 7590
rect 16743 7588 16767 7590
rect 16823 7588 16847 7590
rect 16903 7588 16927 7590
rect 16983 7588 16989 7590
rect 16681 7579 16989 7588
rect 16681 6556 16989 6565
rect 16681 6554 16687 6556
rect 16743 6554 16767 6556
rect 16823 6554 16847 6556
rect 16903 6554 16927 6556
rect 16983 6554 16989 6556
rect 16743 6502 16745 6554
rect 16925 6502 16927 6554
rect 16681 6500 16687 6502
rect 16743 6500 16767 6502
rect 16823 6500 16847 6502
rect 16903 6500 16927 6502
rect 16983 6500 16989 6502
rect 16681 6491 16989 6500
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5778 15332 6054
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3670 13400 3878
rect 14292 3738 14320 4558
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 14476 2922 14504 4558
rect 14568 3126 14596 5170
rect 14715 4924 15023 4933
rect 14715 4922 14721 4924
rect 14777 4922 14801 4924
rect 14857 4922 14881 4924
rect 14937 4922 14961 4924
rect 15017 4922 15023 4924
rect 14777 4870 14779 4922
rect 14959 4870 14961 4922
rect 14715 4868 14721 4870
rect 14777 4868 14801 4870
rect 14857 4868 14881 4870
rect 14937 4868 14961 4870
rect 15017 4868 15023 4870
rect 14715 4859 15023 4868
rect 15212 4826 15240 5714
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 14715 3836 15023 3845
rect 14715 3834 14721 3836
rect 14777 3834 14801 3836
rect 14857 3834 14881 3836
rect 14937 3834 14961 3836
rect 15017 3834 15023 3836
rect 14777 3782 14779 3834
rect 14959 3782 14961 3834
rect 14715 3780 14721 3782
rect 14777 3780 14801 3782
rect 14857 3780 14881 3782
rect 14937 3780 14961 3782
rect 15017 3780 15023 3782
rect 14715 3771 15023 3780
rect 15120 3670 15148 4558
rect 15304 4146 15332 5510
rect 16681 5468 16989 5477
rect 16681 5466 16687 5468
rect 16743 5466 16767 5468
rect 16823 5466 16847 5468
rect 16903 5466 16927 5468
rect 16983 5466 16989 5468
rect 16743 5414 16745 5466
rect 16925 5414 16927 5466
rect 16681 5412 16687 5414
rect 16743 5412 16767 5414
rect 16823 5412 16847 5414
rect 16903 5412 16927 5414
rect 16983 5412 16989 5414
rect 16681 5403 16989 5412
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15488 3194 15516 4082
rect 16040 3534 16068 4422
rect 16316 4146 16344 5102
rect 16681 4380 16989 4389
rect 16681 4378 16687 4380
rect 16743 4378 16767 4380
rect 16823 4378 16847 4380
rect 16903 4378 16927 4380
rect 16983 4378 16989 4380
rect 16743 4326 16745 4378
rect 16925 4326 16927 4378
rect 16681 4324 16687 4326
rect 16743 4324 16767 4326
rect 16823 4324 16847 4326
rect 16903 4324 16927 4326
rect 16983 4324 16989 4326
rect 16681 4315 16989 4324
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12748 2204 13056 2213
rect 12748 2202 12754 2204
rect 12810 2202 12834 2204
rect 12890 2202 12914 2204
rect 12970 2202 12994 2204
rect 13050 2202 13056 2204
rect 12810 2150 12812 2202
rect 12992 2150 12994 2202
rect 12748 2148 12754 2150
rect 12810 2148 12834 2150
rect 12890 2148 12914 2150
rect 12970 2148 12994 2150
rect 13050 2148 13056 2150
rect 12748 2139 13056 2148
rect 13372 800 13400 2858
rect 14568 2446 14596 3062
rect 14715 2748 15023 2757
rect 14715 2746 14721 2748
rect 14777 2746 14801 2748
rect 14857 2746 14881 2748
rect 14937 2746 14961 2748
rect 15017 2746 15023 2748
rect 14777 2694 14779 2746
rect 14959 2694 14961 2746
rect 14715 2692 14721 2694
rect 14777 2692 14801 2694
rect 14857 2692 14881 2694
rect 14937 2692 14961 2694
rect 15017 2692 15023 2694
rect 14715 2683 15023 2692
rect 16224 2582 16252 3470
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16316 3058 16344 3334
rect 16681 3292 16989 3301
rect 16681 3290 16687 3292
rect 16743 3290 16767 3292
rect 16823 3290 16847 3292
rect 16903 3290 16927 3292
rect 16983 3290 16989 3292
rect 16743 3238 16745 3290
rect 16925 3238 16927 3290
rect 16681 3236 16687 3238
rect 16743 3236 16767 3238
rect 16823 3236 16847 3238
rect 16903 3236 16927 3238
rect 16983 3236 16989 3238
rect 16681 3227 16989 3236
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 16316 800 16344 2994
rect 16681 2204 16989 2213
rect 16681 2202 16687 2204
rect 16743 2202 16767 2204
rect 16823 2202 16847 2204
rect 16903 2202 16927 2204
rect 16983 2202 16989 2204
rect 16743 2150 16745 2202
rect 16925 2150 16927 2202
rect 16681 2148 16687 2150
rect 16743 2148 16767 2150
rect 16823 2148 16847 2150
rect 16903 2148 16927 2150
rect 16983 2148 16989 2150
rect 16681 2139 16989 2148
rect 1582 0 1638 800
rect 4526 0 4582 800
rect 7470 0 7526 800
rect 10414 0 10470 800
rect 13358 0 13414 800
rect 16302 0 16358 800
<< via2 >>
rect 2922 15802 2978 15804
rect 3002 15802 3058 15804
rect 3082 15802 3138 15804
rect 3162 15802 3218 15804
rect 2922 15750 2968 15802
rect 2968 15750 2978 15802
rect 3002 15750 3032 15802
rect 3032 15750 3044 15802
rect 3044 15750 3058 15802
rect 3082 15750 3096 15802
rect 3096 15750 3108 15802
rect 3108 15750 3138 15802
rect 3162 15750 3172 15802
rect 3172 15750 3218 15802
rect 2922 15748 2978 15750
rect 3002 15748 3058 15750
rect 3082 15748 3138 15750
rect 3162 15748 3218 15750
rect 6855 15802 6911 15804
rect 6935 15802 6991 15804
rect 7015 15802 7071 15804
rect 7095 15802 7151 15804
rect 6855 15750 6901 15802
rect 6901 15750 6911 15802
rect 6935 15750 6965 15802
rect 6965 15750 6977 15802
rect 6977 15750 6991 15802
rect 7015 15750 7029 15802
rect 7029 15750 7041 15802
rect 7041 15750 7071 15802
rect 7095 15750 7105 15802
rect 7105 15750 7151 15802
rect 6855 15748 6911 15750
rect 6935 15748 6991 15750
rect 7015 15748 7071 15750
rect 7095 15748 7151 15750
rect 10788 15802 10844 15804
rect 10868 15802 10924 15804
rect 10948 15802 11004 15804
rect 11028 15802 11084 15804
rect 10788 15750 10834 15802
rect 10834 15750 10844 15802
rect 10868 15750 10898 15802
rect 10898 15750 10910 15802
rect 10910 15750 10924 15802
rect 10948 15750 10962 15802
rect 10962 15750 10974 15802
rect 10974 15750 11004 15802
rect 11028 15750 11038 15802
rect 11038 15750 11084 15802
rect 10788 15748 10844 15750
rect 10868 15748 10924 15750
rect 10948 15748 11004 15750
rect 11028 15748 11084 15750
rect 14721 15802 14777 15804
rect 14801 15802 14857 15804
rect 14881 15802 14937 15804
rect 14961 15802 15017 15804
rect 14721 15750 14767 15802
rect 14767 15750 14777 15802
rect 14801 15750 14831 15802
rect 14831 15750 14843 15802
rect 14843 15750 14857 15802
rect 14881 15750 14895 15802
rect 14895 15750 14907 15802
rect 14907 15750 14937 15802
rect 14961 15750 14971 15802
rect 14971 15750 15017 15802
rect 14721 15748 14777 15750
rect 14801 15748 14857 15750
rect 14881 15748 14937 15750
rect 14961 15748 15017 15750
rect 2922 14714 2978 14716
rect 3002 14714 3058 14716
rect 3082 14714 3138 14716
rect 3162 14714 3218 14716
rect 2922 14662 2968 14714
rect 2968 14662 2978 14714
rect 3002 14662 3032 14714
rect 3032 14662 3044 14714
rect 3044 14662 3058 14714
rect 3082 14662 3096 14714
rect 3096 14662 3108 14714
rect 3108 14662 3138 14714
rect 3162 14662 3172 14714
rect 3172 14662 3218 14714
rect 2922 14660 2978 14662
rect 3002 14660 3058 14662
rect 3082 14660 3138 14662
rect 3162 14660 3218 14662
rect 2922 13626 2978 13628
rect 3002 13626 3058 13628
rect 3082 13626 3138 13628
rect 3162 13626 3218 13628
rect 2922 13574 2968 13626
rect 2968 13574 2978 13626
rect 3002 13574 3032 13626
rect 3032 13574 3044 13626
rect 3044 13574 3058 13626
rect 3082 13574 3096 13626
rect 3096 13574 3108 13626
rect 3108 13574 3138 13626
rect 3162 13574 3172 13626
rect 3172 13574 3218 13626
rect 2922 13572 2978 13574
rect 3002 13572 3058 13574
rect 3082 13572 3138 13574
rect 3162 13572 3218 13574
rect 2922 12538 2978 12540
rect 3002 12538 3058 12540
rect 3082 12538 3138 12540
rect 3162 12538 3218 12540
rect 2922 12486 2968 12538
rect 2968 12486 2978 12538
rect 3002 12486 3032 12538
rect 3032 12486 3044 12538
rect 3044 12486 3058 12538
rect 3082 12486 3096 12538
rect 3096 12486 3108 12538
rect 3108 12486 3138 12538
rect 3162 12486 3172 12538
rect 3172 12486 3218 12538
rect 2922 12484 2978 12486
rect 3002 12484 3058 12486
rect 3082 12484 3138 12486
rect 3162 12484 3218 12486
rect 2922 11450 2978 11452
rect 3002 11450 3058 11452
rect 3082 11450 3138 11452
rect 3162 11450 3218 11452
rect 2922 11398 2968 11450
rect 2968 11398 2978 11450
rect 3002 11398 3032 11450
rect 3032 11398 3044 11450
rect 3044 11398 3058 11450
rect 3082 11398 3096 11450
rect 3096 11398 3108 11450
rect 3108 11398 3138 11450
rect 3162 11398 3172 11450
rect 3172 11398 3218 11450
rect 2922 11396 2978 11398
rect 3002 11396 3058 11398
rect 3082 11396 3138 11398
rect 3162 11396 3218 11398
rect 2922 10362 2978 10364
rect 3002 10362 3058 10364
rect 3082 10362 3138 10364
rect 3162 10362 3218 10364
rect 2922 10310 2968 10362
rect 2968 10310 2978 10362
rect 3002 10310 3032 10362
rect 3032 10310 3044 10362
rect 3044 10310 3058 10362
rect 3082 10310 3096 10362
rect 3096 10310 3108 10362
rect 3108 10310 3138 10362
rect 3162 10310 3172 10362
rect 3172 10310 3218 10362
rect 2922 10308 2978 10310
rect 3002 10308 3058 10310
rect 3082 10308 3138 10310
rect 3162 10308 3218 10310
rect 2922 9274 2978 9276
rect 3002 9274 3058 9276
rect 3082 9274 3138 9276
rect 3162 9274 3218 9276
rect 2922 9222 2968 9274
rect 2968 9222 2978 9274
rect 3002 9222 3032 9274
rect 3032 9222 3044 9274
rect 3044 9222 3058 9274
rect 3082 9222 3096 9274
rect 3096 9222 3108 9274
rect 3108 9222 3138 9274
rect 3162 9222 3172 9274
rect 3172 9222 3218 9274
rect 2922 9220 2978 9222
rect 3002 9220 3058 9222
rect 3082 9220 3138 9222
rect 3162 9220 3218 9222
rect 2922 8186 2978 8188
rect 3002 8186 3058 8188
rect 3082 8186 3138 8188
rect 3162 8186 3218 8188
rect 2922 8134 2968 8186
rect 2968 8134 2978 8186
rect 3002 8134 3032 8186
rect 3032 8134 3044 8186
rect 3044 8134 3058 8186
rect 3082 8134 3096 8186
rect 3096 8134 3108 8186
rect 3108 8134 3138 8186
rect 3162 8134 3172 8186
rect 3172 8134 3218 8186
rect 2922 8132 2978 8134
rect 3002 8132 3058 8134
rect 3082 8132 3138 8134
rect 3162 8132 3218 8134
rect 2922 7098 2978 7100
rect 3002 7098 3058 7100
rect 3082 7098 3138 7100
rect 3162 7098 3218 7100
rect 2922 7046 2968 7098
rect 2968 7046 2978 7098
rect 3002 7046 3032 7098
rect 3032 7046 3044 7098
rect 3044 7046 3058 7098
rect 3082 7046 3096 7098
rect 3096 7046 3108 7098
rect 3108 7046 3138 7098
rect 3162 7046 3172 7098
rect 3172 7046 3218 7098
rect 2922 7044 2978 7046
rect 3002 7044 3058 7046
rect 3082 7044 3138 7046
rect 3162 7044 3218 7046
rect 2922 6010 2978 6012
rect 3002 6010 3058 6012
rect 3082 6010 3138 6012
rect 3162 6010 3218 6012
rect 2922 5958 2968 6010
rect 2968 5958 2978 6010
rect 3002 5958 3032 6010
rect 3032 5958 3044 6010
rect 3044 5958 3058 6010
rect 3082 5958 3096 6010
rect 3096 5958 3108 6010
rect 3108 5958 3138 6010
rect 3162 5958 3172 6010
rect 3172 5958 3218 6010
rect 2922 5956 2978 5958
rect 3002 5956 3058 5958
rect 3082 5956 3138 5958
rect 3162 5956 3218 5958
rect 4888 15258 4944 15260
rect 4968 15258 5024 15260
rect 5048 15258 5104 15260
rect 5128 15258 5184 15260
rect 4888 15206 4934 15258
rect 4934 15206 4944 15258
rect 4968 15206 4998 15258
rect 4998 15206 5010 15258
rect 5010 15206 5024 15258
rect 5048 15206 5062 15258
rect 5062 15206 5074 15258
rect 5074 15206 5104 15258
rect 5128 15206 5138 15258
rect 5138 15206 5184 15258
rect 4888 15204 4944 15206
rect 4968 15204 5024 15206
rect 5048 15204 5104 15206
rect 5128 15204 5184 15206
rect 8821 15258 8877 15260
rect 8901 15258 8957 15260
rect 8981 15258 9037 15260
rect 9061 15258 9117 15260
rect 8821 15206 8867 15258
rect 8867 15206 8877 15258
rect 8901 15206 8931 15258
rect 8931 15206 8943 15258
rect 8943 15206 8957 15258
rect 8981 15206 8995 15258
rect 8995 15206 9007 15258
rect 9007 15206 9037 15258
rect 9061 15206 9071 15258
rect 9071 15206 9117 15258
rect 8821 15204 8877 15206
rect 8901 15204 8957 15206
rect 8981 15204 9037 15206
rect 9061 15204 9117 15206
rect 6855 14714 6911 14716
rect 6935 14714 6991 14716
rect 7015 14714 7071 14716
rect 7095 14714 7151 14716
rect 6855 14662 6901 14714
rect 6901 14662 6911 14714
rect 6935 14662 6965 14714
rect 6965 14662 6977 14714
rect 6977 14662 6991 14714
rect 7015 14662 7029 14714
rect 7029 14662 7041 14714
rect 7041 14662 7071 14714
rect 7095 14662 7105 14714
rect 7105 14662 7151 14714
rect 6855 14660 6911 14662
rect 6935 14660 6991 14662
rect 7015 14660 7071 14662
rect 7095 14660 7151 14662
rect 4888 14170 4944 14172
rect 4968 14170 5024 14172
rect 5048 14170 5104 14172
rect 5128 14170 5184 14172
rect 4888 14118 4934 14170
rect 4934 14118 4944 14170
rect 4968 14118 4998 14170
rect 4998 14118 5010 14170
rect 5010 14118 5024 14170
rect 5048 14118 5062 14170
rect 5062 14118 5074 14170
rect 5074 14118 5104 14170
rect 5128 14118 5138 14170
rect 5138 14118 5184 14170
rect 4888 14116 4944 14118
rect 4968 14116 5024 14118
rect 5048 14116 5104 14118
rect 5128 14116 5184 14118
rect 8821 14170 8877 14172
rect 8901 14170 8957 14172
rect 8981 14170 9037 14172
rect 9061 14170 9117 14172
rect 8821 14118 8867 14170
rect 8867 14118 8877 14170
rect 8901 14118 8931 14170
rect 8931 14118 8943 14170
rect 8943 14118 8957 14170
rect 8981 14118 8995 14170
rect 8995 14118 9007 14170
rect 9007 14118 9037 14170
rect 9061 14118 9071 14170
rect 9071 14118 9117 14170
rect 8821 14116 8877 14118
rect 8901 14116 8957 14118
rect 8981 14116 9037 14118
rect 9061 14116 9117 14118
rect 6855 13626 6911 13628
rect 6935 13626 6991 13628
rect 7015 13626 7071 13628
rect 7095 13626 7151 13628
rect 6855 13574 6901 13626
rect 6901 13574 6911 13626
rect 6935 13574 6965 13626
rect 6965 13574 6977 13626
rect 6977 13574 6991 13626
rect 7015 13574 7029 13626
rect 7029 13574 7041 13626
rect 7041 13574 7071 13626
rect 7095 13574 7105 13626
rect 7105 13574 7151 13626
rect 6855 13572 6911 13574
rect 6935 13572 6991 13574
rect 7015 13572 7071 13574
rect 7095 13572 7151 13574
rect 4888 13082 4944 13084
rect 4968 13082 5024 13084
rect 5048 13082 5104 13084
rect 5128 13082 5184 13084
rect 4888 13030 4934 13082
rect 4934 13030 4944 13082
rect 4968 13030 4998 13082
rect 4998 13030 5010 13082
rect 5010 13030 5024 13082
rect 5048 13030 5062 13082
rect 5062 13030 5074 13082
rect 5074 13030 5104 13082
rect 5128 13030 5138 13082
rect 5138 13030 5184 13082
rect 4888 13028 4944 13030
rect 4968 13028 5024 13030
rect 5048 13028 5104 13030
rect 5128 13028 5184 13030
rect 8821 13082 8877 13084
rect 8901 13082 8957 13084
rect 8981 13082 9037 13084
rect 9061 13082 9117 13084
rect 8821 13030 8867 13082
rect 8867 13030 8877 13082
rect 8901 13030 8931 13082
rect 8931 13030 8943 13082
rect 8943 13030 8957 13082
rect 8981 13030 8995 13082
rect 8995 13030 9007 13082
rect 9007 13030 9037 13082
rect 9061 13030 9071 13082
rect 9071 13030 9117 13082
rect 8821 13028 8877 13030
rect 8901 13028 8957 13030
rect 8981 13028 9037 13030
rect 9061 13028 9117 13030
rect 6855 12538 6911 12540
rect 6935 12538 6991 12540
rect 7015 12538 7071 12540
rect 7095 12538 7151 12540
rect 6855 12486 6901 12538
rect 6901 12486 6911 12538
rect 6935 12486 6965 12538
rect 6965 12486 6977 12538
rect 6977 12486 6991 12538
rect 7015 12486 7029 12538
rect 7029 12486 7041 12538
rect 7041 12486 7071 12538
rect 7095 12486 7105 12538
rect 7105 12486 7151 12538
rect 6855 12484 6911 12486
rect 6935 12484 6991 12486
rect 7015 12484 7071 12486
rect 7095 12484 7151 12486
rect 4888 11994 4944 11996
rect 4968 11994 5024 11996
rect 5048 11994 5104 11996
rect 5128 11994 5184 11996
rect 4888 11942 4934 11994
rect 4934 11942 4944 11994
rect 4968 11942 4998 11994
rect 4998 11942 5010 11994
rect 5010 11942 5024 11994
rect 5048 11942 5062 11994
rect 5062 11942 5074 11994
rect 5074 11942 5104 11994
rect 5128 11942 5138 11994
rect 5138 11942 5184 11994
rect 4888 11940 4944 11942
rect 4968 11940 5024 11942
rect 5048 11940 5104 11942
rect 5128 11940 5184 11942
rect 8821 11994 8877 11996
rect 8901 11994 8957 11996
rect 8981 11994 9037 11996
rect 9061 11994 9117 11996
rect 8821 11942 8867 11994
rect 8867 11942 8877 11994
rect 8901 11942 8931 11994
rect 8931 11942 8943 11994
rect 8943 11942 8957 11994
rect 8981 11942 8995 11994
rect 8995 11942 9007 11994
rect 9007 11942 9037 11994
rect 9061 11942 9071 11994
rect 9071 11942 9117 11994
rect 8821 11940 8877 11942
rect 8901 11940 8957 11942
rect 8981 11940 9037 11942
rect 9061 11940 9117 11942
rect 6855 11450 6911 11452
rect 6935 11450 6991 11452
rect 7015 11450 7071 11452
rect 7095 11450 7151 11452
rect 6855 11398 6901 11450
rect 6901 11398 6911 11450
rect 6935 11398 6965 11450
rect 6965 11398 6977 11450
rect 6977 11398 6991 11450
rect 7015 11398 7029 11450
rect 7029 11398 7041 11450
rect 7041 11398 7071 11450
rect 7095 11398 7105 11450
rect 7105 11398 7151 11450
rect 6855 11396 6911 11398
rect 6935 11396 6991 11398
rect 7015 11396 7071 11398
rect 7095 11396 7151 11398
rect 4888 10906 4944 10908
rect 4968 10906 5024 10908
rect 5048 10906 5104 10908
rect 5128 10906 5184 10908
rect 4888 10854 4934 10906
rect 4934 10854 4944 10906
rect 4968 10854 4998 10906
rect 4998 10854 5010 10906
rect 5010 10854 5024 10906
rect 5048 10854 5062 10906
rect 5062 10854 5074 10906
rect 5074 10854 5104 10906
rect 5128 10854 5138 10906
rect 5138 10854 5184 10906
rect 4888 10852 4944 10854
rect 4968 10852 5024 10854
rect 5048 10852 5104 10854
rect 5128 10852 5184 10854
rect 8821 10906 8877 10908
rect 8901 10906 8957 10908
rect 8981 10906 9037 10908
rect 9061 10906 9117 10908
rect 8821 10854 8867 10906
rect 8867 10854 8877 10906
rect 8901 10854 8931 10906
rect 8931 10854 8943 10906
rect 8943 10854 8957 10906
rect 8981 10854 8995 10906
rect 8995 10854 9007 10906
rect 9007 10854 9037 10906
rect 9061 10854 9071 10906
rect 9071 10854 9117 10906
rect 8821 10852 8877 10854
rect 8901 10852 8957 10854
rect 8981 10852 9037 10854
rect 9061 10852 9117 10854
rect 6855 10362 6911 10364
rect 6935 10362 6991 10364
rect 7015 10362 7071 10364
rect 7095 10362 7151 10364
rect 6855 10310 6901 10362
rect 6901 10310 6911 10362
rect 6935 10310 6965 10362
rect 6965 10310 6977 10362
rect 6977 10310 6991 10362
rect 7015 10310 7029 10362
rect 7029 10310 7041 10362
rect 7041 10310 7071 10362
rect 7095 10310 7105 10362
rect 7105 10310 7151 10362
rect 6855 10308 6911 10310
rect 6935 10308 6991 10310
rect 7015 10308 7071 10310
rect 7095 10308 7151 10310
rect 4888 9818 4944 9820
rect 4968 9818 5024 9820
rect 5048 9818 5104 9820
rect 5128 9818 5184 9820
rect 4888 9766 4934 9818
rect 4934 9766 4944 9818
rect 4968 9766 4998 9818
rect 4998 9766 5010 9818
rect 5010 9766 5024 9818
rect 5048 9766 5062 9818
rect 5062 9766 5074 9818
rect 5074 9766 5104 9818
rect 5128 9766 5138 9818
rect 5138 9766 5184 9818
rect 4888 9764 4944 9766
rect 4968 9764 5024 9766
rect 5048 9764 5104 9766
rect 5128 9764 5184 9766
rect 8821 9818 8877 9820
rect 8901 9818 8957 9820
rect 8981 9818 9037 9820
rect 9061 9818 9117 9820
rect 8821 9766 8867 9818
rect 8867 9766 8877 9818
rect 8901 9766 8931 9818
rect 8931 9766 8943 9818
rect 8943 9766 8957 9818
rect 8981 9766 8995 9818
rect 8995 9766 9007 9818
rect 9007 9766 9037 9818
rect 9061 9766 9071 9818
rect 9071 9766 9117 9818
rect 8821 9764 8877 9766
rect 8901 9764 8957 9766
rect 8981 9764 9037 9766
rect 9061 9764 9117 9766
rect 6855 9274 6911 9276
rect 6935 9274 6991 9276
rect 7015 9274 7071 9276
rect 7095 9274 7151 9276
rect 6855 9222 6901 9274
rect 6901 9222 6911 9274
rect 6935 9222 6965 9274
rect 6965 9222 6977 9274
rect 6977 9222 6991 9274
rect 7015 9222 7029 9274
rect 7029 9222 7041 9274
rect 7041 9222 7071 9274
rect 7095 9222 7105 9274
rect 7105 9222 7151 9274
rect 6855 9220 6911 9222
rect 6935 9220 6991 9222
rect 7015 9220 7071 9222
rect 7095 9220 7151 9222
rect 4888 8730 4944 8732
rect 4968 8730 5024 8732
rect 5048 8730 5104 8732
rect 5128 8730 5184 8732
rect 4888 8678 4934 8730
rect 4934 8678 4944 8730
rect 4968 8678 4998 8730
rect 4998 8678 5010 8730
rect 5010 8678 5024 8730
rect 5048 8678 5062 8730
rect 5062 8678 5074 8730
rect 5074 8678 5104 8730
rect 5128 8678 5138 8730
rect 5138 8678 5184 8730
rect 4888 8676 4944 8678
rect 4968 8676 5024 8678
rect 5048 8676 5104 8678
rect 5128 8676 5184 8678
rect 8821 8730 8877 8732
rect 8901 8730 8957 8732
rect 8981 8730 9037 8732
rect 9061 8730 9117 8732
rect 8821 8678 8867 8730
rect 8867 8678 8877 8730
rect 8901 8678 8931 8730
rect 8931 8678 8943 8730
rect 8943 8678 8957 8730
rect 8981 8678 8995 8730
rect 8995 8678 9007 8730
rect 9007 8678 9037 8730
rect 9061 8678 9071 8730
rect 9071 8678 9117 8730
rect 8821 8676 8877 8678
rect 8901 8676 8957 8678
rect 8981 8676 9037 8678
rect 9061 8676 9117 8678
rect 6855 8186 6911 8188
rect 6935 8186 6991 8188
rect 7015 8186 7071 8188
rect 7095 8186 7151 8188
rect 6855 8134 6901 8186
rect 6901 8134 6911 8186
rect 6935 8134 6965 8186
rect 6965 8134 6977 8186
rect 6977 8134 6991 8186
rect 7015 8134 7029 8186
rect 7029 8134 7041 8186
rect 7041 8134 7071 8186
rect 7095 8134 7105 8186
rect 7105 8134 7151 8186
rect 6855 8132 6911 8134
rect 6935 8132 6991 8134
rect 7015 8132 7071 8134
rect 7095 8132 7151 8134
rect 4888 7642 4944 7644
rect 4968 7642 5024 7644
rect 5048 7642 5104 7644
rect 5128 7642 5184 7644
rect 4888 7590 4934 7642
rect 4934 7590 4944 7642
rect 4968 7590 4998 7642
rect 4998 7590 5010 7642
rect 5010 7590 5024 7642
rect 5048 7590 5062 7642
rect 5062 7590 5074 7642
rect 5074 7590 5104 7642
rect 5128 7590 5138 7642
rect 5138 7590 5184 7642
rect 4888 7588 4944 7590
rect 4968 7588 5024 7590
rect 5048 7588 5104 7590
rect 5128 7588 5184 7590
rect 8821 7642 8877 7644
rect 8901 7642 8957 7644
rect 8981 7642 9037 7644
rect 9061 7642 9117 7644
rect 8821 7590 8867 7642
rect 8867 7590 8877 7642
rect 8901 7590 8931 7642
rect 8931 7590 8943 7642
rect 8943 7590 8957 7642
rect 8981 7590 8995 7642
rect 8995 7590 9007 7642
rect 9007 7590 9037 7642
rect 9061 7590 9071 7642
rect 9071 7590 9117 7642
rect 8821 7588 8877 7590
rect 8901 7588 8957 7590
rect 8981 7588 9037 7590
rect 9061 7588 9117 7590
rect 6855 7098 6911 7100
rect 6935 7098 6991 7100
rect 7015 7098 7071 7100
rect 7095 7098 7151 7100
rect 6855 7046 6901 7098
rect 6901 7046 6911 7098
rect 6935 7046 6965 7098
rect 6965 7046 6977 7098
rect 6977 7046 6991 7098
rect 7015 7046 7029 7098
rect 7029 7046 7041 7098
rect 7041 7046 7071 7098
rect 7095 7046 7105 7098
rect 7105 7046 7151 7098
rect 6855 7044 6911 7046
rect 6935 7044 6991 7046
rect 7015 7044 7071 7046
rect 7095 7044 7151 7046
rect 4888 6554 4944 6556
rect 4968 6554 5024 6556
rect 5048 6554 5104 6556
rect 5128 6554 5184 6556
rect 4888 6502 4934 6554
rect 4934 6502 4944 6554
rect 4968 6502 4998 6554
rect 4998 6502 5010 6554
rect 5010 6502 5024 6554
rect 5048 6502 5062 6554
rect 5062 6502 5074 6554
rect 5074 6502 5104 6554
rect 5128 6502 5138 6554
rect 5138 6502 5184 6554
rect 4888 6500 4944 6502
rect 4968 6500 5024 6502
rect 5048 6500 5104 6502
rect 5128 6500 5184 6502
rect 8821 6554 8877 6556
rect 8901 6554 8957 6556
rect 8981 6554 9037 6556
rect 9061 6554 9117 6556
rect 8821 6502 8867 6554
rect 8867 6502 8877 6554
rect 8901 6502 8931 6554
rect 8931 6502 8943 6554
rect 8943 6502 8957 6554
rect 8981 6502 8995 6554
rect 8995 6502 9007 6554
rect 9007 6502 9037 6554
rect 9061 6502 9071 6554
rect 9071 6502 9117 6554
rect 8821 6500 8877 6502
rect 8901 6500 8957 6502
rect 8981 6500 9037 6502
rect 9061 6500 9117 6502
rect 6855 6010 6911 6012
rect 6935 6010 6991 6012
rect 7015 6010 7071 6012
rect 7095 6010 7151 6012
rect 6855 5958 6901 6010
rect 6901 5958 6911 6010
rect 6935 5958 6965 6010
rect 6965 5958 6977 6010
rect 6977 5958 6991 6010
rect 7015 5958 7029 6010
rect 7029 5958 7041 6010
rect 7041 5958 7071 6010
rect 7095 5958 7105 6010
rect 7105 5958 7151 6010
rect 6855 5956 6911 5958
rect 6935 5956 6991 5958
rect 7015 5956 7071 5958
rect 7095 5956 7151 5958
rect 4888 5466 4944 5468
rect 4968 5466 5024 5468
rect 5048 5466 5104 5468
rect 5128 5466 5184 5468
rect 4888 5414 4934 5466
rect 4934 5414 4944 5466
rect 4968 5414 4998 5466
rect 4998 5414 5010 5466
rect 5010 5414 5024 5466
rect 5048 5414 5062 5466
rect 5062 5414 5074 5466
rect 5074 5414 5104 5466
rect 5128 5414 5138 5466
rect 5138 5414 5184 5466
rect 4888 5412 4944 5414
rect 4968 5412 5024 5414
rect 5048 5412 5104 5414
rect 5128 5412 5184 5414
rect 8821 5466 8877 5468
rect 8901 5466 8957 5468
rect 8981 5466 9037 5468
rect 9061 5466 9117 5468
rect 8821 5414 8867 5466
rect 8867 5414 8877 5466
rect 8901 5414 8931 5466
rect 8931 5414 8943 5466
rect 8943 5414 8957 5466
rect 8981 5414 8995 5466
rect 8995 5414 9007 5466
rect 9007 5414 9037 5466
rect 9061 5414 9071 5466
rect 9071 5414 9117 5466
rect 8821 5412 8877 5414
rect 8901 5412 8957 5414
rect 8981 5412 9037 5414
rect 9061 5412 9117 5414
rect 2922 4922 2978 4924
rect 3002 4922 3058 4924
rect 3082 4922 3138 4924
rect 3162 4922 3218 4924
rect 2922 4870 2968 4922
rect 2968 4870 2978 4922
rect 3002 4870 3032 4922
rect 3032 4870 3044 4922
rect 3044 4870 3058 4922
rect 3082 4870 3096 4922
rect 3096 4870 3108 4922
rect 3108 4870 3138 4922
rect 3162 4870 3172 4922
rect 3172 4870 3218 4922
rect 2922 4868 2978 4870
rect 3002 4868 3058 4870
rect 3082 4868 3138 4870
rect 3162 4868 3218 4870
rect 6855 4922 6911 4924
rect 6935 4922 6991 4924
rect 7015 4922 7071 4924
rect 7095 4922 7151 4924
rect 6855 4870 6901 4922
rect 6901 4870 6911 4922
rect 6935 4870 6965 4922
rect 6965 4870 6977 4922
rect 6977 4870 6991 4922
rect 7015 4870 7029 4922
rect 7029 4870 7041 4922
rect 7041 4870 7071 4922
rect 7095 4870 7105 4922
rect 7105 4870 7151 4922
rect 6855 4868 6911 4870
rect 6935 4868 6991 4870
rect 7015 4868 7071 4870
rect 7095 4868 7151 4870
rect 4888 4378 4944 4380
rect 4968 4378 5024 4380
rect 5048 4378 5104 4380
rect 5128 4378 5184 4380
rect 4888 4326 4934 4378
rect 4934 4326 4944 4378
rect 4968 4326 4998 4378
rect 4998 4326 5010 4378
rect 5010 4326 5024 4378
rect 5048 4326 5062 4378
rect 5062 4326 5074 4378
rect 5074 4326 5104 4378
rect 5128 4326 5138 4378
rect 5138 4326 5184 4378
rect 4888 4324 4944 4326
rect 4968 4324 5024 4326
rect 5048 4324 5104 4326
rect 5128 4324 5184 4326
rect 8821 4378 8877 4380
rect 8901 4378 8957 4380
rect 8981 4378 9037 4380
rect 9061 4378 9117 4380
rect 8821 4326 8867 4378
rect 8867 4326 8877 4378
rect 8901 4326 8931 4378
rect 8931 4326 8943 4378
rect 8943 4326 8957 4378
rect 8981 4326 8995 4378
rect 8995 4326 9007 4378
rect 9007 4326 9037 4378
rect 9061 4326 9071 4378
rect 9071 4326 9117 4378
rect 8821 4324 8877 4326
rect 8901 4324 8957 4326
rect 8981 4324 9037 4326
rect 9061 4324 9117 4326
rect 12754 15258 12810 15260
rect 12834 15258 12890 15260
rect 12914 15258 12970 15260
rect 12994 15258 13050 15260
rect 12754 15206 12800 15258
rect 12800 15206 12810 15258
rect 12834 15206 12864 15258
rect 12864 15206 12876 15258
rect 12876 15206 12890 15258
rect 12914 15206 12928 15258
rect 12928 15206 12940 15258
rect 12940 15206 12970 15258
rect 12994 15206 13004 15258
rect 13004 15206 13050 15258
rect 12754 15204 12810 15206
rect 12834 15204 12890 15206
rect 12914 15204 12970 15206
rect 12994 15204 13050 15206
rect 10788 14714 10844 14716
rect 10868 14714 10924 14716
rect 10948 14714 11004 14716
rect 11028 14714 11084 14716
rect 10788 14662 10834 14714
rect 10834 14662 10844 14714
rect 10868 14662 10898 14714
rect 10898 14662 10910 14714
rect 10910 14662 10924 14714
rect 10948 14662 10962 14714
rect 10962 14662 10974 14714
rect 10974 14662 11004 14714
rect 11028 14662 11038 14714
rect 11038 14662 11084 14714
rect 10788 14660 10844 14662
rect 10868 14660 10924 14662
rect 10948 14660 11004 14662
rect 11028 14660 11084 14662
rect 12754 14170 12810 14172
rect 12834 14170 12890 14172
rect 12914 14170 12970 14172
rect 12994 14170 13050 14172
rect 12754 14118 12800 14170
rect 12800 14118 12810 14170
rect 12834 14118 12864 14170
rect 12864 14118 12876 14170
rect 12876 14118 12890 14170
rect 12914 14118 12928 14170
rect 12928 14118 12940 14170
rect 12940 14118 12970 14170
rect 12994 14118 13004 14170
rect 13004 14118 13050 14170
rect 12754 14116 12810 14118
rect 12834 14116 12890 14118
rect 12914 14116 12970 14118
rect 12994 14116 13050 14118
rect 10788 13626 10844 13628
rect 10868 13626 10924 13628
rect 10948 13626 11004 13628
rect 11028 13626 11084 13628
rect 10788 13574 10834 13626
rect 10834 13574 10844 13626
rect 10868 13574 10898 13626
rect 10898 13574 10910 13626
rect 10910 13574 10924 13626
rect 10948 13574 10962 13626
rect 10962 13574 10974 13626
rect 10974 13574 11004 13626
rect 11028 13574 11038 13626
rect 11038 13574 11084 13626
rect 10788 13572 10844 13574
rect 10868 13572 10924 13574
rect 10948 13572 11004 13574
rect 11028 13572 11084 13574
rect 12754 13082 12810 13084
rect 12834 13082 12890 13084
rect 12914 13082 12970 13084
rect 12994 13082 13050 13084
rect 12754 13030 12800 13082
rect 12800 13030 12810 13082
rect 12834 13030 12864 13082
rect 12864 13030 12876 13082
rect 12876 13030 12890 13082
rect 12914 13030 12928 13082
rect 12928 13030 12940 13082
rect 12940 13030 12970 13082
rect 12994 13030 13004 13082
rect 13004 13030 13050 13082
rect 12754 13028 12810 13030
rect 12834 13028 12890 13030
rect 12914 13028 12970 13030
rect 12994 13028 13050 13030
rect 10788 12538 10844 12540
rect 10868 12538 10924 12540
rect 10948 12538 11004 12540
rect 11028 12538 11084 12540
rect 10788 12486 10834 12538
rect 10834 12486 10844 12538
rect 10868 12486 10898 12538
rect 10898 12486 10910 12538
rect 10910 12486 10924 12538
rect 10948 12486 10962 12538
rect 10962 12486 10974 12538
rect 10974 12486 11004 12538
rect 11028 12486 11038 12538
rect 11038 12486 11084 12538
rect 10788 12484 10844 12486
rect 10868 12484 10924 12486
rect 10948 12484 11004 12486
rect 11028 12484 11084 12486
rect 12754 11994 12810 11996
rect 12834 11994 12890 11996
rect 12914 11994 12970 11996
rect 12994 11994 13050 11996
rect 12754 11942 12800 11994
rect 12800 11942 12810 11994
rect 12834 11942 12864 11994
rect 12864 11942 12876 11994
rect 12876 11942 12890 11994
rect 12914 11942 12928 11994
rect 12928 11942 12940 11994
rect 12940 11942 12970 11994
rect 12994 11942 13004 11994
rect 13004 11942 13050 11994
rect 12754 11940 12810 11942
rect 12834 11940 12890 11942
rect 12914 11940 12970 11942
rect 12994 11940 13050 11942
rect 10788 11450 10844 11452
rect 10868 11450 10924 11452
rect 10948 11450 11004 11452
rect 11028 11450 11084 11452
rect 10788 11398 10834 11450
rect 10834 11398 10844 11450
rect 10868 11398 10898 11450
rect 10898 11398 10910 11450
rect 10910 11398 10924 11450
rect 10948 11398 10962 11450
rect 10962 11398 10974 11450
rect 10974 11398 11004 11450
rect 11028 11398 11038 11450
rect 11038 11398 11084 11450
rect 10788 11396 10844 11398
rect 10868 11396 10924 11398
rect 10948 11396 11004 11398
rect 11028 11396 11084 11398
rect 12754 10906 12810 10908
rect 12834 10906 12890 10908
rect 12914 10906 12970 10908
rect 12994 10906 13050 10908
rect 12754 10854 12800 10906
rect 12800 10854 12810 10906
rect 12834 10854 12864 10906
rect 12864 10854 12876 10906
rect 12876 10854 12890 10906
rect 12914 10854 12928 10906
rect 12928 10854 12940 10906
rect 12940 10854 12970 10906
rect 12994 10854 13004 10906
rect 13004 10854 13050 10906
rect 12754 10852 12810 10854
rect 12834 10852 12890 10854
rect 12914 10852 12970 10854
rect 12994 10852 13050 10854
rect 10788 10362 10844 10364
rect 10868 10362 10924 10364
rect 10948 10362 11004 10364
rect 11028 10362 11084 10364
rect 10788 10310 10834 10362
rect 10834 10310 10844 10362
rect 10868 10310 10898 10362
rect 10898 10310 10910 10362
rect 10910 10310 10924 10362
rect 10948 10310 10962 10362
rect 10962 10310 10974 10362
rect 10974 10310 11004 10362
rect 11028 10310 11038 10362
rect 11038 10310 11084 10362
rect 10788 10308 10844 10310
rect 10868 10308 10924 10310
rect 10948 10308 11004 10310
rect 11028 10308 11084 10310
rect 12754 9818 12810 9820
rect 12834 9818 12890 9820
rect 12914 9818 12970 9820
rect 12994 9818 13050 9820
rect 12754 9766 12800 9818
rect 12800 9766 12810 9818
rect 12834 9766 12864 9818
rect 12864 9766 12876 9818
rect 12876 9766 12890 9818
rect 12914 9766 12928 9818
rect 12928 9766 12940 9818
rect 12940 9766 12970 9818
rect 12994 9766 13004 9818
rect 13004 9766 13050 9818
rect 12754 9764 12810 9766
rect 12834 9764 12890 9766
rect 12914 9764 12970 9766
rect 12994 9764 13050 9766
rect 10788 9274 10844 9276
rect 10868 9274 10924 9276
rect 10948 9274 11004 9276
rect 11028 9274 11084 9276
rect 10788 9222 10834 9274
rect 10834 9222 10844 9274
rect 10868 9222 10898 9274
rect 10898 9222 10910 9274
rect 10910 9222 10924 9274
rect 10948 9222 10962 9274
rect 10962 9222 10974 9274
rect 10974 9222 11004 9274
rect 11028 9222 11038 9274
rect 11038 9222 11084 9274
rect 10788 9220 10844 9222
rect 10868 9220 10924 9222
rect 10948 9220 11004 9222
rect 11028 9220 11084 9222
rect 12754 8730 12810 8732
rect 12834 8730 12890 8732
rect 12914 8730 12970 8732
rect 12994 8730 13050 8732
rect 12754 8678 12800 8730
rect 12800 8678 12810 8730
rect 12834 8678 12864 8730
rect 12864 8678 12876 8730
rect 12876 8678 12890 8730
rect 12914 8678 12928 8730
rect 12928 8678 12940 8730
rect 12940 8678 12970 8730
rect 12994 8678 13004 8730
rect 13004 8678 13050 8730
rect 12754 8676 12810 8678
rect 12834 8676 12890 8678
rect 12914 8676 12970 8678
rect 12994 8676 13050 8678
rect 10788 8186 10844 8188
rect 10868 8186 10924 8188
rect 10948 8186 11004 8188
rect 11028 8186 11084 8188
rect 10788 8134 10834 8186
rect 10834 8134 10844 8186
rect 10868 8134 10898 8186
rect 10898 8134 10910 8186
rect 10910 8134 10924 8186
rect 10948 8134 10962 8186
rect 10962 8134 10974 8186
rect 10974 8134 11004 8186
rect 11028 8134 11038 8186
rect 11038 8134 11084 8186
rect 10788 8132 10844 8134
rect 10868 8132 10924 8134
rect 10948 8132 11004 8134
rect 11028 8132 11084 8134
rect 12754 7642 12810 7644
rect 12834 7642 12890 7644
rect 12914 7642 12970 7644
rect 12994 7642 13050 7644
rect 12754 7590 12800 7642
rect 12800 7590 12810 7642
rect 12834 7590 12864 7642
rect 12864 7590 12876 7642
rect 12876 7590 12890 7642
rect 12914 7590 12928 7642
rect 12928 7590 12940 7642
rect 12940 7590 12970 7642
rect 12994 7590 13004 7642
rect 13004 7590 13050 7642
rect 12754 7588 12810 7590
rect 12834 7588 12890 7590
rect 12914 7588 12970 7590
rect 12994 7588 13050 7590
rect 10788 7098 10844 7100
rect 10868 7098 10924 7100
rect 10948 7098 11004 7100
rect 11028 7098 11084 7100
rect 10788 7046 10834 7098
rect 10834 7046 10844 7098
rect 10868 7046 10898 7098
rect 10898 7046 10910 7098
rect 10910 7046 10924 7098
rect 10948 7046 10962 7098
rect 10962 7046 10974 7098
rect 10974 7046 11004 7098
rect 11028 7046 11038 7098
rect 11038 7046 11084 7098
rect 10788 7044 10844 7046
rect 10868 7044 10924 7046
rect 10948 7044 11004 7046
rect 11028 7044 11084 7046
rect 10788 6010 10844 6012
rect 10868 6010 10924 6012
rect 10948 6010 11004 6012
rect 11028 6010 11084 6012
rect 10788 5958 10834 6010
rect 10834 5958 10844 6010
rect 10868 5958 10898 6010
rect 10898 5958 10910 6010
rect 10910 5958 10924 6010
rect 10948 5958 10962 6010
rect 10962 5958 10974 6010
rect 10974 5958 11004 6010
rect 11028 5958 11038 6010
rect 11038 5958 11084 6010
rect 10788 5956 10844 5958
rect 10868 5956 10924 5958
rect 10948 5956 11004 5958
rect 11028 5956 11084 5958
rect 12754 6554 12810 6556
rect 12834 6554 12890 6556
rect 12914 6554 12970 6556
rect 12994 6554 13050 6556
rect 12754 6502 12800 6554
rect 12800 6502 12810 6554
rect 12834 6502 12864 6554
rect 12864 6502 12876 6554
rect 12876 6502 12890 6554
rect 12914 6502 12928 6554
rect 12928 6502 12940 6554
rect 12940 6502 12970 6554
rect 12994 6502 13004 6554
rect 13004 6502 13050 6554
rect 12754 6500 12810 6502
rect 12834 6500 12890 6502
rect 12914 6500 12970 6502
rect 12994 6500 13050 6502
rect 10788 4922 10844 4924
rect 10868 4922 10924 4924
rect 10948 4922 11004 4924
rect 11028 4922 11084 4924
rect 10788 4870 10834 4922
rect 10834 4870 10844 4922
rect 10868 4870 10898 4922
rect 10898 4870 10910 4922
rect 10910 4870 10924 4922
rect 10948 4870 10962 4922
rect 10962 4870 10974 4922
rect 10974 4870 11004 4922
rect 11028 4870 11038 4922
rect 11038 4870 11084 4922
rect 10788 4868 10844 4870
rect 10868 4868 10924 4870
rect 10948 4868 11004 4870
rect 11028 4868 11084 4870
rect 2922 3834 2978 3836
rect 3002 3834 3058 3836
rect 3082 3834 3138 3836
rect 3162 3834 3218 3836
rect 2922 3782 2968 3834
rect 2968 3782 2978 3834
rect 3002 3782 3032 3834
rect 3032 3782 3044 3834
rect 3044 3782 3058 3834
rect 3082 3782 3096 3834
rect 3096 3782 3108 3834
rect 3108 3782 3138 3834
rect 3162 3782 3172 3834
rect 3172 3782 3218 3834
rect 2922 3780 2978 3782
rect 3002 3780 3058 3782
rect 3082 3780 3138 3782
rect 3162 3780 3218 3782
rect 6855 3834 6911 3836
rect 6935 3834 6991 3836
rect 7015 3834 7071 3836
rect 7095 3834 7151 3836
rect 6855 3782 6901 3834
rect 6901 3782 6911 3834
rect 6935 3782 6965 3834
rect 6965 3782 6977 3834
rect 6977 3782 6991 3834
rect 7015 3782 7029 3834
rect 7029 3782 7041 3834
rect 7041 3782 7071 3834
rect 7095 3782 7105 3834
rect 7105 3782 7151 3834
rect 6855 3780 6911 3782
rect 6935 3780 6991 3782
rect 7015 3780 7071 3782
rect 7095 3780 7151 3782
rect 4888 3290 4944 3292
rect 4968 3290 5024 3292
rect 5048 3290 5104 3292
rect 5128 3290 5184 3292
rect 4888 3238 4934 3290
rect 4934 3238 4944 3290
rect 4968 3238 4998 3290
rect 4998 3238 5010 3290
rect 5010 3238 5024 3290
rect 5048 3238 5062 3290
rect 5062 3238 5074 3290
rect 5074 3238 5104 3290
rect 5128 3238 5138 3290
rect 5138 3238 5184 3290
rect 4888 3236 4944 3238
rect 4968 3236 5024 3238
rect 5048 3236 5104 3238
rect 5128 3236 5184 3238
rect 8821 3290 8877 3292
rect 8901 3290 8957 3292
rect 8981 3290 9037 3292
rect 9061 3290 9117 3292
rect 8821 3238 8867 3290
rect 8867 3238 8877 3290
rect 8901 3238 8931 3290
rect 8931 3238 8943 3290
rect 8943 3238 8957 3290
rect 8981 3238 8995 3290
rect 8995 3238 9007 3290
rect 9007 3238 9037 3290
rect 9061 3238 9071 3290
rect 9071 3238 9117 3290
rect 8821 3236 8877 3238
rect 8901 3236 8957 3238
rect 8981 3236 9037 3238
rect 9061 3236 9117 3238
rect 2922 2746 2978 2748
rect 3002 2746 3058 2748
rect 3082 2746 3138 2748
rect 3162 2746 3218 2748
rect 2922 2694 2968 2746
rect 2968 2694 2978 2746
rect 3002 2694 3032 2746
rect 3032 2694 3044 2746
rect 3044 2694 3058 2746
rect 3082 2694 3096 2746
rect 3096 2694 3108 2746
rect 3108 2694 3138 2746
rect 3162 2694 3172 2746
rect 3172 2694 3218 2746
rect 2922 2692 2978 2694
rect 3002 2692 3058 2694
rect 3082 2692 3138 2694
rect 3162 2692 3218 2694
rect 6855 2746 6911 2748
rect 6935 2746 6991 2748
rect 7015 2746 7071 2748
rect 7095 2746 7151 2748
rect 6855 2694 6901 2746
rect 6901 2694 6911 2746
rect 6935 2694 6965 2746
rect 6965 2694 6977 2746
rect 6977 2694 6991 2746
rect 7015 2694 7029 2746
rect 7029 2694 7041 2746
rect 7041 2694 7071 2746
rect 7095 2694 7105 2746
rect 7105 2694 7151 2746
rect 6855 2692 6911 2694
rect 6935 2692 6991 2694
rect 7015 2692 7071 2694
rect 7095 2692 7151 2694
rect 4888 2202 4944 2204
rect 4968 2202 5024 2204
rect 5048 2202 5104 2204
rect 5128 2202 5184 2204
rect 4888 2150 4934 2202
rect 4934 2150 4944 2202
rect 4968 2150 4998 2202
rect 4998 2150 5010 2202
rect 5010 2150 5024 2202
rect 5048 2150 5062 2202
rect 5062 2150 5074 2202
rect 5074 2150 5104 2202
rect 5128 2150 5138 2202
rect 5138 2150 5184 2202
rect 4888 2148 4944 2150
rect 4968 2148 5024 2150
rect 5048 2148 5104 2150
rect 5128 2148 5184 2150
rect 10788 3834 10844 3836
rect 10868 3834 10924 3836
rect 10948 3834 11004 3836
rect 11028 3834 11084 3836
rect 10788 3782 10834 3834
rect 10834 3782 10844 3834
rect 10868 3782 10898 3834
rect 10898 3782 10910 3834
rect 10910 3782 10924 3834
rect 10948 3782 10962 3834
rect 10962 3782 10974 3834
rect 10974 3782 11004 3834
rect 11028 3782 11038 3834
rect 11038 3782 11084 3834
rect 10788 3780 10844 3782
rect 10868 3780 10924 3782
rect 10948 3780 11004 3782
rect 11028 3780 11084 3782
rect 10788 2746 10844 2748
rect 10868 2746 10924 2748
rect 10948 2746 11004 2748
rect 11028 2746 11084 2748
rect 10788 2694 10834 2746
rect 10834 2694 10844 2746
rect 10868 2694 10898 2746
rect 10898 2694 10910 2746
rect 10910 2694 10924 2746
rect 10948 2694 10962 2746
rect 10962 2694 10974 2746
rect 10974 2694 11004 2746
rect 11028 2694 11038 2746
rect 11038 2694 11084 2746
rect 10788 2692 10844 2694
rect 10868 2692 10924 2694
rect 10948 2692 11004 2694
rect 11028 2692 11084 2694
rect 8821 2202 8877 2204
rect 8901 2202 8957 2204
rect 8981 2202 9037 2204
rect 9061 2202 9117 2204
rect 8821 2150 8867 2202
rect 8867 2150 8877 2202
rect 8901 2150 8931 2202
rect 8931 2150 8943 2202
rect 8943 2150 8957 2202
rect 8981 2150 8995 2202
rect 8995 2150 9007 2202
rect 9007 2150 9037 2202
rect 9061 2150 9071 2202
rect 9071 2150 9117 2202
rect 8821 2148 8877 2150
rect 8901 2148 8957 2150
rect 8981 2148 9037 2150
rect 9061 2148 9117 2150
rect 12754 5466 12810 5468
rect 12834 5466 12890 5468
rect 12914 5466 12970 5468
rect 12994 5466 13050 5468
rect 12754 5414 12800 5466
rect 12800 5414 12810 5466
rect 12834 5414 12864 5466
rect 12864 5414 12876 5466
rect 12876 5414 12890 5466
rect 12914 5414 12928 5466
rect 12928 5414 12940 5466
rect 12940 5414 12970 5466
rect 12994 5414 13004 5466
rect 13004 5414 13050 5466
rect 12754 5412 12810 5414
rect 12834 5412 12890 5414
rect 12914 5412 12970 5414
rect 12994 5412 13050 5414
rect 12754 4378 12810 4380
rect 12834 4378 12890 4380
rect 12914 4378 12970 4380
rect 12994 4378 13050 4380
rect 12754 4326 12800 4378
rect 12800 4326 12810 4378
rect 12834 4326 12864 4378
rect 12864 4326 12876 4378
rect 12876 4326 12890 4378
rect 12914 4326 12928 4378
rect 12928 4326 12940 4378
rect 12940 4326 12970 4378
rect 12994 4326 13004 4378
rect 13004 4326 13050 4378
rect 12754 4324 12810 4326
rect 12834 4324 12890 4326
rect 12914 4324 12970 4326
rect 12994 4324 13050 4326
rect 12754 3290 12810 3292
rect 12834 3290 12890 3292
rect 12914 3290 12970 3292
rect 12994 3290 13050 3292
rect 12754 3238 12800 3290
rect 12800 3238 12810 3290
rect 12834 3238 12864 3290
rect 12864 3238 12876 3290
rect 12876 3238 12890 3290
rect 12914 3238 12928 3290
rect 12928 3238 12940 3290
rect 12940 3238 12970 3290
rect 12994 3238 13004 3290
rect 13004 3238 13050 3290
rect 12754 3236 12810 3238
rect 12834 3236 12890 3238
rect 12914 3236 12970 3238
rect 12994 3236 13050 3238
rect 14721 14714 14777 14716
rect 14801 14714 14857 14716
rect 14881 14714 14937 14716
rect 14961 14714 15017 14716
rect 14721 14662 14767 14714
rect 14767 14662 14777 14714
rect 14801 14662 14831 14714
rect 14831 14662 14843 14714
rect 14843 14662 14857 14714
rect 14881 14662 14895 14714
rect 14895 14662 14907 14714
rect 14907 14662 14937 14714
rect 14961 14662 14971 14714
rect 14971 14662 15017 14714
rect 14721 14660 14777 14662
rect 14801 14660 14857 14662
rect 14881 14660 14937 14662
rect 14961 14660 15017 14662
rect 14721 13626 14777 13628
rect 14801 13626 14857 13628
rect 14881 13626 14937 13628
rect 14961 13626 15017 13628
rect 14721 13574 14767 13626
rect 14767 13574 14777 13626
rect 14801 13574 14831 13626
rect 14831 13574 14843 13626
rect 14843 13574 14857 13626
rect 14881 13574 14895 13626
rect 14895 13574 14907 13626
rect 14907 13574 14937 13626
rect 14961 13574 14971 13626
rect 14971 13574 15017 13626
rect 14721 13572 14777 13574
rect 14801 13572 14857 13574
rect 14881 13572 14937 13574
rect 14961 13572 15017 13574
rect 14721 12538 14777 12540
rect 14801 12538 14857 12540
rect 14881 12538 14937 12540
rect 14961 12538 15017 12540
rect 14721 12486 14767 12538
rect 14767 12486 14777 12538
rect 14801 12486 14831 12538
rect 14831 12486 14843 12538
rect 14843 12486 14857 12538
rect 14881 12486 14895 12538
rect 14895 12486 14907 12538
rect 14907 12486 14937 12538
rect 14961 12486 14971 12538
rect 14971 12486 15017 12538
rect 14721 12484 14777 12486
rect 14801 12484 14857 12486
rect 14881 12484 14937 12486
rect 14961 12484 15017 12486
rect 14721 11450 14777 11452
rect 14801 11450 14857 11452
rect 14881 11450 14937 11452
rect 14961 11450 15017 11452
rect 14721 11398 14767 11450
rect 14767 11398 14777 11450
rect 14801 11398 14831 11450
rect 14831 11398 14843 11450
rect 14843 11398 14857 11450
rect 14881 11398 14895 11450
rect 14895 11398 14907 11450
rect 14907 11398 14937 11450
rect 14961 11398 14971 11450
rect 14971 11398 15017 11450
rect 14721 11396 14777 11398
rect 14801 11396 14857 11398
rect 14881 11396 14937 11398
rect 14961 11396 15017 11398
rect 14721 10362 14777 10364
rect 14801 10362 14857 10364
rect 14881 10362 14937 10364
rect 14961 10362 15017 10364
rect 14721 10310 14767 10362
rect 14767 10310 14777 10362
rect 14801 10310 14831 10362
rect 14831 10310 14843 10362
rect 14843 10310 14857 10362
rect 14881 10310 14895 10362
rect 14895 10310 14907 10362
rect 14907 10310 14937 10362
rect 14961 10310 14971 10362
rect 14971 10310 15017 10362
rect 14721 10308 14777 10310
rect 14801 10308 14857 10310
rect 14881 10308 14937 10310
rect 14961 10308 15017 10310
rect 14721 9274 14777 9276
rect 14801 9274 14857 9276
rect 14881 9274 14937 9276
rect 14961 9274 15017 9276
rect 14721 9222 14767 9274
rect 14767 9222 14777 9274
rect 14801 9222 14831 9274
rect 14831 9222 14843 9274
rect 14843 9222 14857 9274
rect 14881 9222 14895 9274
rect 14895 9222 14907 9274
rect 14907 9222 14937 9274
rect 14961 9222 14971 9274
rect 14971 9222 15017 9274
rect 14721 9220 14777 9222
rect 14801 9220 14857 9222
rect 14881 9220 14937 9222
rect 14961 9220 15017 9222
rect 14721 8186 14777 8188
rect 14801 8186 14857 8188
rect 14881 8186 14937 8188
rect 14961 8186 15017 8188
rect 14721 8134 14767 8186
rect 14767 8134 14777 8186
rect 14801 8134 14831 8186
rect 14831 8134 14843 8186
rect 14843 8134 14857 8186
rect 14881 8134 14895 8186
rect 14895 8134 14907 8186
rect 14907 8134 14937 8186
rect 14961 8134 14971 8186
rect 14971 8134 15017 8186
rect 14721 8132 14777 8134
rect 14801 8132 14857 8134
rect 14881 8132 14937 8134
rect 14961 8132 15017 8134
rect 14721 7098 14777 7100
rect 14801 7098 14857 7100
rect 14881 7098 14937 7100
rect 14961 7098 15017 7100
rect 14721 7046 14767 7098
rect 14767 7046 14777 7098
rect 14801 7046 14831 7098
rect 14831 7046 14843 7098
rect 14843 7046 14857 7098
rect 14881 7046 14895 7098
rect 14895 7046 14907 7098
rect 14907 7046 14937 7098
rect 14961 7046 14971 7098
rect 14971 7046 15017 7098
rect 14721 7044 14777 7046
rect 14801 7044 14857 7046
rect 14881 7044 14937 7046
rect 14961 7044 15017 7046
rect 14721 6010 14777 6012
rect 14801 6010 14857 6012
rect 14881 6010 14937 6012
rect 14961 6010 15017 6012
rect 14721 5958 14767 6010
rect 14767 5958 14777 6010
rect 14801 5958 14831 6010
rect 14831 5958 14843 6010
rect 14843 5958 14857 6010
rect 14881 5958 14895 6010
rect 14895 5958 14907 6010
rect 14907 5958 14937 6010
rect 14961 5958 14971 6010
rect 14971 5958 15017 6010
rect 14721 5956 14777 5958
rect 14801 5956 14857 5958
rect 14881 5956 14937 5958
rect 14961 5956 15017 5958
rect 16687 15258 16743 15260
rect 16767 15258 16823 15260
rect 16847 15258 16903 15260
rect 16927 15258 16983 15260
rect 16687 15206 16733 15258
rect 16733 15206 16743 15258
rect 16767 15206 16797 15258
rect 16797 15206 16809 15258
rect 16809 15206 16823 15258
rect 16847 15206 16861 15258
rect 16861 15206 16873 15258
rect 16873 15206 16903 15258
rect 16927 15206 16937 15258
rect 16937 15206 16983 15258
rect 16687 15204 16743 15206
rect 16767 15204 16823 15206
rect 16847 15204 16903 15206
rect 16927 15204 16983 15206
rect 16687 14170 16743 14172
rect 16767 14170 16823 14172
rect 16847 14170 16903 14172
rect 16927 14170 16983 14172
rect 16687 14118 16733 14170
rect 16733 14118 16743 14170
rect 16767 14118 16797 14170
rect 16797 14118 16809 14170
rect 16809 14118 16823 14170
rect 16847 14118 16861 14170
rect 16861 14118 16873 14170
rect 16873 14118 16903 14170
rect 16927 14118 16937 14170
rect 16937 14118 16983 14170
rect 16687 14116 16743 14118
rect 16767 14116 16823 14118
rect 16847 14116 16903 14118
rect 16927 14116 16983 14118
rect 16687 13082 16743 13084
rect 16767 13082 16823 13084
rect 16847 13082 16903 13084
rect 16927 13082 16983 13084
rect 16687 13030 16733 13082
rect 16733 13030 16743 13082
rect 16767 13030 16797 13082
rect 16797 13030 16809 13082
rect 16809 13030 16823 13082
rect 16847 13030 16861 13082
rect 16861 13030 16873 13082
rect 16873 13030 16903 13082
rect 16927 13030 16937 13082
rect 16937 13030 16983 13082
rect 16687 13028 16743 13030
rect 16767 13028 16823 13030
rect 16847 13028 16903 13030
rect 16927 13028 16983 13030
rect 16687 11994 16743 11996
rect 16767 11994 16823 11996
rect 16847 11994 16903 11996
rect 16927 11994 16983 11996
rect 16687 11942 16733 11994
rect 16733 11942 16743 11994
rect 16767 11942 16797 11994
rect 16797 11942 16809 11994
rect 16809 11942 16823 11994
rect 16847 11942 16861 11994
rect 16861 11942 16873 11994
rect 16873 11942 16903 11994
rect 16927 11942 16937 11994
rect 16937 11942 16983 11994
rect 16687 11940 16743 11942
rect 16767 11940 16823 11942
rect 16847 11940 16903 11942
rect 16927 11940 16983 11942
rect 16687 10906 16743 10908
rect 16767 10906 16823 10908
rect 16847 10906 16903 10908
rect 16927 10906 16983 10908
rect 16687 10854 16733 10906
rect 16733 10854 16743 10906
rect 16767 10854 16797 10906
rect 16797 10854 16809 10906
rect 16809 10854 16823 10906
rect 16847 10854 16861 10906
rect 16861 10854 16873 10906
rect 16873 10854 16903 10906
rect 16927 10854 16937 10906
rect 16937 10854 16983 10906
rect 16687 10852 16743 10854
rect 16767 10852 16823 10854
rect 16847 10852 16903 10854
rect 16927 10852 16983 10854
rect 16687 9818 16743 9820
rect 16767 9818 16823 9820
rect 16847 9818 16903 9820
rect 16927 9818 16983 9820
rect 16687 9766 16733 9818
rect 16733 9766 16743 9818
rect 16767 9766 16797 9818
rect 16797 9766 16809 9818
rect 16809 9766 16823 9818
rect 16847 9766 16861 9818
rect 16861 9766 16873 9818
rect 16873 9766 16903 9818
rect 16927 9766 16937 9818
rect 16937 9766 16983 9818
rect 16687 9764 16743 9766
rect 16767 9764 16823 9766
rect 16847 9764 16903 9766
rect 16927 9764 16983 9766
rect 16687 8730 16743 8732
rect 16767 8730 16823 8732
rect 16847 8730 16903 8732
rect 16927 8730 16983 8732
rect 16687 8678 16733 8730
rect 16733 8678 16743 8730
rect 16767 8678 16797 8730
rect 16797 8678 16809 8730
rect 16809 8678 16823 8730
rect 16847 8678 16861 8730
rect 16861 8678 16873 8730
rect 16873 8678 16903 8730
rect 16927 8678 16937 8730
rect 16937 8678 16983 8730
rect 16687 8676 16743 8678
rect 16767 8676 16823 8678
rect 16847 8676 16903 8678
rect 16927 8676 16983 8678
rect 16687 7642 16743 7644
rect 16767 7642 16823 7644
rect 16847 7642 16903 7644
rect 16927 7642 16983 7644
rect 16687 7590 16733 7642
rect 16733 7590 16743 7642
rect 16767 7590 16797 7642
rect 16797 7590 16809 7642
rect 16809 7590 16823 7642
rect 16847 7590 16861 7642
rect 16861 7590 16873 7642
rect 16873 7590 16903 7642
rect 16927 7590 16937 7642
rect 16937 7590 16983 7642
rect 16687 7588 16743 7590
rect 16767 7588 16823 7590
rect 16847 7588 16903 7590
rect 16927 7588 16983 7590
rect 16687 6554 16743 6556
rect 16767 6554 16823 6556
rect 16847 6554 16903 6556
rect 16927 6554 16983 6556
rect 16687 6502 16733 6554
rect 16733 6502 16743 6554
rect 16767 6502 16797 6554
rect 16797 6502 16809 6554
rect 16809 6502 16823 6554
rect 16847 6502 16861 6554
rect 16861 6502 16873 6554
rect 16873 6502 16903 6554
rect 16927 6502 16937 6554
rect 16937 6502 16983 6554
rect 16687 6500 16743 6502
rect 16767 6500 16823 6502
rect 16847 6500 16903 6502
rect 16927 6500 16983 6502
rect 14721 4922 14777 4924
rect 14801 4922 14857 4924
rect 14881 4922 14937 4924
rect 14961 4922 15017 4924
rect 14721 4870 14767 4922
rect 14767 4870 14777 4922
rect 14801 4870 14831 4922
rect 14831 4870 14843 4922
rect 14843 4870 14857 4922
rect 14881 4870 14895 4922
rect 14895 4870 14907 4922
rect 14907 4870 14937 4922
rect 14961 4870 14971 4922
rect 14971 4870 15017 4922
rect 14721 4868 14777 4870
rect 14801 4868 14857 4870
rect 14881 4868 14937 4870
rect 14961 4868 15017 4870
rect 14721 3834 14777 3836
rect 14801 3834 14857 3836
rect 14881 3834 14937 3836
rect 14961 3834 15017 3836
rect 14721 3782 14767 3834
rect 14767 3782 14777 3834
rect 14801 3782 14831 3834
rect 14831 3782 14843 3834
rect 14843 3782 14857 3834
rect 14881 3782 14895 3834
rect 14895 3782 14907 3834
rect 14907 3782 14937 3834
rect 14961 3782 14971 3834
rect 14971 3782 15017 3834
rect 14721 3780 14777 3782
rect 14801 3780 14857 3782
rect 14881 3780 14937 3782
rect 14961 3780 15017 3782
rect 16687 5466 16743 5468
rect 16767 5466 16823 5468
rect 16847 5466 16903 5468
rect 16927 5466 16983 5468
rect 16687 5414 16733 5466
rect 16733 5414 16743 5466
rect 16767 5414 16797 5466
rect 16797 5414 16809 5466
rect 16809 5414 16823 5466
rect 16847 5414 16861 5466
rect 16861 5414 16873 5466
rect 16873 5414 16903 5466
rect 16927 5414 16937 5466
rect 16937 5414 16983 5466
rect 16687 5412 16743 5414
rect 16767 5412 16823 5414
rect 16847 5412 16903 5414
rect 16927 5412 16983 5414
rect 16687 4378 16743 4380
rect 16767 4378 16823 4380
rect 16847 4378 16903 4380
rect 16927 4378 16983 4380
rect 16687 4326 16733 4378
rect 16733 4326 16743 4378
rect 16767 4326 16797 4378
rect 16797 4326 16809 4378
rect 16809 4326 16823 4378
rect 16847 4326 16861 4378
rect 16861 4326 16873 4378
rect 16873 4326 16903 4378
rect 16927 4326 16937 4378
rect 16937 4326 16983 4378
rect 16687 4324 16743 4326
rect 16767 4324 16823 4326
rect 16847 4324 16903 4326
rect 16927 4324 16983 4326
rect 12754 2202 12810 2204
rect 12834 2202 12890 2204
rect 12914 2202 12970 2204
rect 12994 2202 13050 2204
rect 12754 2150 12800 2202
rect 12800 2150 12810 2202
rect 12834 2150 12864 2202
rect 12864 2150 12876 2202
rect 12876 2150 12890 2202
rect 12914 2150 12928 2202
rect 12928 2150 12940 2202
rect 12940 2150 12970 2202
rect 12994 2150 13004 2202
rect 13004 2150 13050 2202
rect 12754 2148 12810 2150
rect 12834 2148 12890 2150
rect 12914 2148 12970 2150
rect 12994 2148 13050 2150
rect 14721 2746 14777 2748
rect 14801 2746 14857 2748
rect 14881 2746 14937 2748
rect 14961 2746 15017 2748
rect 14721 2694 14767 2746
rect 14767 2694 14777 2746
rect 14801 2694 14831 2746
rect 14831 2694 14843 2746
rect 14843 2694 14857 2746
rect 14881 2694 14895 2746
rect 14895 2694 14907 2746
rect 14907 2694 14937 2746
rect 14961 2694 14971 2746
rect 14971 2694 15017 2746
rect 14721 2692 14777 2694
rect 14801 2692 14857 2694
rect 14881 2692 14937 2694
rect 14961 2692 15017 2694
rect 16687 3290 16743 3292
rect 16767 3290 16823 3292
rect 16847 3290 16903 3292
rect 16927 3290 16983 3292
rect 16687 3238 16733 3290
rect 16733 3238 16743 3290
rect 16767 3238 16797 3290
rect 16797 3238 16809 3290
rect 16809 3238 16823 3290
rect 16847 3238 16861 3290
rect 16861 3238 16873 3290
rect 16873 3238 16903 3290
rect 16927 3238 16937 3290
rect 16937 3238 16983 3290
rect 16687 3236 16743 3238
rect 16767 3236 16823 3238
rect 16847 3236 16903 3238
rect 16927 3236 16983 3238
rect 16687 2202 16743 2204
rect 16767 2202 16823 2204
rect 16847 2202 16903 2204
rect 16927 2202 16983 2204
rect 16687 2150 16733 2202
rect 16733 2150 16743 2202
rect 16767 2150 16797 2202
rect 16797 2150 16809 2202
rect 16809 2150 16823 2202
rect 16847 2150 16861 2202
rect 16861 2150 16873 2202
rect 16873 2150 16903 2202
rect 16927 2150 16937 2202
rect 16937 2150 16983 2202
rect 16687 2148 16743 2150
rect 16767 2148 16823 2150
rect 16847 2148 16903 2150
rect 16927 2148 16983 2150
<< metal3 >>
rect 2912 15808 3228 15809
rect 2912 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3228 15808
rect 2912 15743 3228 15744
rect 6845 15808 7161 15809
rect 6845 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7161 15808
rect 6845 15743 7161 15744
rect 10778 15808 11094 15809
rect 10778 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11094 15808
rect 10778 15743 11094 15744
rect 14711 15808 15027 15809
rect 14711 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15027 15808
rect 14711 15743 15027 15744
rect 4878 15264 5194 15265
rect 4878 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5194 15264
rect 4878 15199 5194 15200
rect 8811 15264 9127 15265
rect 8811 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9127 15264
rect 8811 15199 9127 15200
rect 12744 15264 13060 15265
rect 12744 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13060 15264
rect 12744 15199 13060 15200
rect 16677 15264 16993 15265
rect 16677 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16993 15264
rect 16677 15199 16993 15200
rect 2912 14720 3228 14721
rect 2912 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3228 14720
rect 2912 14655 3228 14656
rect 6845 14720 7161 14721
rect 6845 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7161 14720
rect 6845 14655 7161 14656
rect 10778 14720 11094 14721
rect 10778 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11094 14720
rect 10778 14655 11094 14656
rect 14711 14720 15027 14721
rect 14711 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15027 14720
rect 14711 14655 15027 14656
rect 4878 14176 5194 14177
rect 4878 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5194 14176
rect 4878 14111 5194 14112
rect 8811 14176 9127 14177
rect 8811 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9127 14176
rect 8811 14111 9127 14112
rect 12744 14176 13060 14177
rect 12744 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13060 14176
rect 12744 14111 13060 14112
rect 16677 14176 16993 14177
rect 16677 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16993 14176
rect 16677 14111 16993 14112
rect 2912 13632 3228 13633
rect 2912 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3228 13632
rect 2912 13567 3228 13568
rect 6845 13632 7161 13633
rect 6845 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7161 13632
rect 6845 13567 7161 13568
rect 10778 13632 11094 13633
rect 10778 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11094 13632
rect 10778 13567 11094 13568
rect 14711 13632 15027 13633
rect 14711 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15027 13632
rect 14711 13567 15027 13568
rect 4878 13088 5194 13089
rect 4878 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5194 13088
rect 4878 13023 5194 13024
rect 8811 13088 9127 13089
rect 8811 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9127 13088
rect 8811 13023 9127 13024
rect 12744 13088 13060 13089
rect 12744 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13060 13088
rect 12744 13023 13060 13024
rect 16677 13088 16993 13089
rect 16677 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16993 13088
rect 16677 13023 16993 13024
rect 2912 12544 3228 12545
rect 2912 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3228 12544
rect 2912 12479 3228 12480
rect 6845 12544 7161 12545
rect 6845 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7161 12544
rect 6845 12479 7161 12480
rect 10778 12544 11094 12545
rect 10778 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11094 12544
rect 10778 12479 11094 12480
rect 14711 12544 15027 12545
rect 14711 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15027 12544
rect 14711 12479 15027 12480
rect 4878 12000 5194 12001
rect 4878 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5194 12000
rect 4878 11935 5194 11936
rect 8811 12000 9127 12001
rect 8811 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9127 12000
rect 8811 11935 9127 11936
rect 12744 12000 13060 12001
rect 12744 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13060 12000
rect 12744 11935 13060 11936
rect 16677 12000 16993 12001
rect 16677 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16993 12000
rect 16677 11935 16993 11936
rect 2912 11456 3228 11457
rect 2912 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3228 11456
rect 2912 11391 3228 11392
rect 6845 11456 7161 11457
rect 6845 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7161 11456
rect 6845 11391 7161 11392
rect 10778 11456 11094 11457
rect 10778 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11094 11456
rect 10778 11391 11094 11392
rect 14711 11456 15027 11457
rect 14711 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15027 11456
rect 14711 11391 15027 11392
rect 4878 10912 5194 10913
rect 4878 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5194 10912
rect 4878 10847 5194 10848
rect 8811 10912 9127 10913
rect 8811 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9127 10912
rect 8811 10847 9127 10848
rect 12744 10912 13060 10913
rect 12744 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13060 10912
rect 12744 10847 13060 10848
rect 16677 10912 16993 10913
rect 16677 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16993 10912
rect 16677 10847 16993 10848
rect 2912 10368 3228 10369
rect 2912 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3228 10368
rect 2912 10303 3228 10304
rect 6845 10368 7161 10369
rect 6845 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7161 10368
rect 6845 10303 7161 10304
rect 10778 10368 11094 10369
rect 10778 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11094 10368
rect 10778 10303 11094 10304
rect 14711 10368 15027 10369
rect 14711 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15027 10368
rect 14711 10303 15027 10304
rect 4878 9824 5194 9825
rect 4878 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5194 9824
rect 4878 9759 5194 9760
rect 8811 9824 9127 9825
rect 8811 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9127 9824
rect 8811 9759 9127 9760
rect 12744 9824 13060 9825
rect 12744 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13060 9824
rect 12744 9759 13060 9760
rect 16677 9824 16993 9825
rect 16677 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16993 9824
rect 16677 9759 16993 9760
rect 2912 9280 3228 9281
rect 2912 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3228 9280
rect 2912 9215 3228 9216
rect 6845 9280 7161 9281
rect 6845 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7161 9280
rect 6845 9215 7161 9216
rect 10778 9280 11094 9281
rect 10778 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11094 9280
rect 10778 9215 11094 9216
rect 14711 9280 15027 9281
rect 14711 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15027 9280
rect 14711 9215 15027 9216
rect 4878 8736 5194 8737
rect 4878 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5194 8736
rect 4878 8671 5194 8672
rect 8811 8736 9127 8737
rect 8811 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9127 8736
rect 8811 8671 9127 8672
rect 12744 8736 13060 8737
rect 12744 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13060 8736
rect 12744 8671 13060 8672
rect 16677 8736 16993 8737
rect 16677 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16993 8736
rect 16677 8671 16993 8672
rect 2912 8192 3228 8193
rect 2912 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3228 8192
rect 2912 8127 3228 8128
rect 6845 8192 7161 8193
rect 6845 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7161 8192
rect 6845 8127 7161 8128
rect 10778 8192 11094 8193
rect 10778 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11094 8192
rect 10778 8127 11094 8128
rect 14711 8192 15027 8193
rect 14711 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15027 8192
rect 14711 8127 15027 8128
rect 4878 7648 5194 7649
rect 4878 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5194 7648
rect 4878 7583 5194 7584
rect 8811 7648 9127 7649
rect 8811 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9127 7648
rect 8811 7583 9127 7584
rect 12744 7648 13060 7649
rect 12744 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13060 7648
rect 12744 7583 13060 7584
rect 16677 7648 16993 7649
rect 16677 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16993 7648
rect 16677 7583 16993 7584
rect 2912 7104 3228 7105
rect 2912 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3228 7104
rect 2912 7039 3228 7040
rect 6845 7104 7161 7105
rect 6845 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7161 7104
rect 6845 7039 7161 7040
rect 10778 7104 11094 7105
rect 10778 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11094 7104
rect 10778 7039 11094 7040
rect 14711 7104 15027 7105
rect 14711 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15027 7104
rect 14711 7039 15027 7040
rect 4878 6560 5194 6561
rect 4878 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5194 6560
rect 4878 6495 5194 6496
rect 8811 6560 9127 6561
rect 8811 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9127 6560
rect 8811 6495 9127 6496
rect 12744 6560 13060 6561
rect 12744 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13060 6560
rect 12744 6495 13060 6496
rect 16677 6560 16993 6561
rect 16677 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16993 6560
rect 16677 6495 16993 6496
rect 2912 6016 3228 6017
rect 2912 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3228 6016
rect 2912 5951 3228 5952
rect 6845 6016 7161 6017
rect 6845 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7161 6016
rect 6845 5951 7161 5952
rect 10778 6016 11094 6017
rect 10778 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11094 6016
rect 10778 5951 11094 5952
rect 14711 6016 15027 6017
rect 14711 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15027 6016
rect 14711 5951 15027 5952
rect 4878 5472 5194 5473
rect 4878 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5194 5472
rect 4878 5407 5194 5408
rect 8811 5472 9127 5473
rect 8811 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9127 5472
rect 8811 5407 9127 5408
rect 12744 5472 13060 5473
rect 12744 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13060 5472
rect 12744 5407 13060 5408
rect 16677 5472 16993 5473
rect 16677 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16993 5472
rect 16677 5407 16993 5408
rect 2912 4928 3228 4929
rect 2912 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3228 4928
rect 2912 4863 3228 4864
rect 6845 4928 7161 4929
rect 6845 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7161 4928
rect 6845 4863 7161 4864
rect 10778 4928 11094 4929
rect 10778 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11094 4928
rect 10778 4863 11094 4864
rect 14711 4928 15027 4929
rect 14711 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15027 4928
rect 14711 4863 15027 4864
rect 4878 4384 5194 4385
rect 4878 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5194 4384
rect 4878 4319 5194 4320
rect 8811 4384 9127 4385
rect 8811 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9127 4384
rect 8811 4319 9127 4320
rect 12744 4384 13060 4385
rect 12744 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13060 4384
rect 12744 4319 13060 4320
rect 16677 4384 16993 4385
rect 16677 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16993 4384
rect 16677 4319 16993 4320
rect 2912 3840 3228 3841
rect 2912 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3228 3840
rect 2912 3775 3228 3776
rect 6845 3840 7161 3841
rect 6845 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7161 3840
rect 6845 3775 7161 3776
rect 10778 3840 11094 3841
rect 10778 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11094 3840
rect 10778 3775 11094 3776
rect 14711 3840 15027 3841
rect 14711 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15027 3840
rect 14711 3775 15027 3776
rect 4878 3296 5194 3297
rect 4878 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5194 3296
rect 4878 3231 5194 3232
rect 8811 3296 9127 3297
rect 8811 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9127 3296
rect 8811 3231 9127 3232
rect 12744 3296 13060 3297
rect 12744 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13060 3296
rect 12744 3231 13060 3232
rect 16677 3296 16993 3297
rect 16677 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16993 3296
rect 16677 3231 16993 3232
rect 2912 2752 3228 2753
rect 2912 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3228 2752
rect 2912 2687 3228 2688
rect 6845 2752 7161 2753
rect 6845 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7161 2752
rect 6845 2687 7161 2688
rect 10778 2752 11094 2753
rect 10778 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11094 2752
rect 10778 2687 11094 2688
rect 14711 2752 15027 2753
rect 14711 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15027 2752
rect 14711 2687 15027 2688
rect 4878 2208 5194 2209
rect 4878 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5194 2208
rect 4878 2143 5194 2144
rect 8811 2208 9127 2209
rect 8811 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9127 2208
rect 8811 2143 9127 2144
rect 12744 2208 13060 2209
rect 12744 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13060 2208
rect 12744 2143 13060 2144
rect 16677 2208 16993 2209
rect 16677 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16993 2208
rect 16677 2143 16993 2144
<< via3 >>
rect 2918 15804 2982 15808
rect 2918 15748 2922 15804
rect 2922 15748 2978 15804
rect 2978 15748 2982 15804
rect 2918 15744 2982 15748
rect 2998 15804 3062 15808
rect 2998 15748 3002 15804
rect 3002 15748 3058 15804
rect 3058 15748 3062 15804
rect 2998 15744 3062 15748
rect 3078 15804 3142 15808
rect 3078 15748 3082 15804
rect 3082 15748 3138 15804
rect 3138 15748 3142 15804
rect 3078 15744 3142 15748
rect 3158 15804 3222 15808
rect 3158 15748 3162 15804
rect 3162 15748 3218 15804
rect 3218 15748 3222 15804
rect 3158 15744 3222 15748
rect 6851 15804 6915 15808
rect 6851 15748 6855 15804
rect 6855 15748 6911 15804
rect 6911 15748 6915 15804
rect 6851 15744 6915 15748
rect 6931 15804 6995 15808
rect 6931 15748 6935 15804
rect 6935 15748 6991 15804
rect 6991 15748 6995 15804
rect 6931 15744 6995 15748
rect 7011 15804 7075 15808
rect 7011 15748 7015 15804
rect 7015 15748 7071 15804
rect 7071 15748 7075 15804
rect 7011 15744 7075 15748
rect 7091 15804 7155 15808
rect 7091 15748 7095 15804
rect 7095 15748 7151 15804
rect 7151 15748 7155 15804
rect 7091 15744 7155 15748
rect 10784 15804 10848 15808
rect 10784 15748 10788 15804
rect 10788 15748 10844 15804
rect 10844 15748 10848 15804
rect 10784 15744 10848 15748
rect 10864 15804 10928 15808
rect 10864 15748 10868 15804
rect 10868 15748 10924 15804
rect 10924 15748 10928 15804
rect 10864 15744 10928 15748
rect 10944 15804 11008 15808
rect 10944 15748 10948 15804
rect 10948 15748 11004 15804
rect 11004 15748 11008 15804
rect 10944 15744 11008 15748
rect 11024 15804 11088 15808
rect 11024 15748 11028 15804
rect 11028 15748 11084 15804
rect 11084 15748 11088 15804
rect 11024 15744 11088 15748
rect 14717 15804 14781 15808
rect 14717 15748 14721 15804
rect 14721 15748 14777 15804
rect 14777 15748 14781 15804
rect 14717 15744 14781 15748
rect 14797 15804 14861 15808
rect 14797 15748 14801 15804
rect 14801 15748 14857 15804
rect 14857 15748 14861 15804
rect 14797 15744 14861 15748
rect 14877 15804 14941 15808
rect 14877 15748 14881 15804
rect 14881 15748 14937 15804
rect 14937 15748 14941 15804
rect 14877 15744 14941 15748
rect 14957 15804 15021 15808
rect 14957 15748 14961 15804
rect 14961 15748 15017 15804
rect 15017 15748 15021 15804
rect 14957 15744 15021 15748
rect 4884 15260 4948 15264
rect 4884 15204 4888 15260
rect 4888 15204 4944 15260
rect 4944 15204 4948 15260
rect 4884 15200 4948 15204
rect 4964 15260 5028 15264
rect 4964 15204 4968 15260
rect 4968 15204 5024 15260
rect 5024 15204 5028 15260
rect 4964 15200 5028 15204
rect 5044 15260 5108 15264
rect 5044 15204 5048 15260
rect 5048 15204 5104 15260
rect 5104 15204 5108 15260
rect 5044 15200 5108 15204
rect 5124 15260 5188 15264
rect 5124 15204 5128 15260
rect 5128 15204 5184 15260
rect 5184 15204 5188 15260
rect 5124 15200 5188 15204
rect 8817 15260 8881 15264
rect 8817 15204 8821 15260
rect 8821 15204 8877 15260
rect 8877 15204 8881 15260
rect 8817 15200 8881 15204
rect 8897 15260 8961 15264
rect 8897 15204 8901 15260
rect 8901 15204 8957 15260
rect 8957 15204 8961 15260
rect 8897 15200 8961 15204
rect 8977 15260 9041 15264
rect 8977 15204 8981 15260
rect 8981 15204 9037 15260
rect 9037 15204 9041 15260
rect 8977 15200 9041 15204
rect 9057 15260 9121 15264
rect 9057 15204 9061 15260
rect 9061 15204 9117 15260
rect 9117 15204 9121 15260
rect 9057 15200 9121 15204
rect 12750 15260 12814 15264
rect 12750 15204 12754 15260
rect 12754 15204 12810 15260
rect 12810 15204 12814 15260
rect 12750 15200 12814 15204
rect 12830 15260 12894 15264
rect 12830 15204 12834 15260
rect 12834 15204 12890 15260
rect 12890 15204 12894 15260
rect 12830 15200 12894 15204
rect 12910 15260 12974 15264
rect 12910 15204 12914 15260
rect 12914 15204 12970 15260
rect 12970 15204 12974 15260
rect 12910 15200 12974 15204
rect 12990 15260 13054 15264
rect 12990 15204 12994 15260
rect 12994 15204 13050 15260
rect 13050 15204 13054 15260
rect 12990 15200 13054 15204
rect 16683 15260 16747 15264
rect 16683 15204 16687 15260
rect 16687 15204 16743 15260
rect 16743 15204 16747 15260
rect 16683 15200 16747 15204
rect 16763 15260 16827 15264
rect 16763 15204 16767 15260
rect 16767 15204 16823 15260
rect 16823 15204 16827 15260
rect 16763 15200 16827 15204
rect 16843 15260 16907 15264
rect 16843 15204 16847 15260
rect 16847 15204 16903 15260
rect 16903 15204 16907 15260
rect 16843 15200 16907 15204
rect 16923 15260 16987 15264
rect 16923 15204 16927 15260
rect 16927 15204 16983 15260
rect 16983 15204 16987 15260
rect 16923 15200 16987 15204
rect 2918 14716 2982 14720
rect 2918 14660 2922 14716
rect 2922 14660 2978 14716
rect 2978 14660 2982 14716
rect 2918 14656 2982 14660
rect 2998 14716 3062 14720
rect 2998 14660 3002 14716
rect 3002 14660 3058 14716
rect 3058 14660 3062 14716
rect 2998 14656 3062 14660
rect 3078 14716 3142 14720
rect 3078 14660 3082 14716
rect 3082 14660 3138 14716
rect 3138 14660 3142 14716
rect 3078 14656 3142 14660
rect 3158 14716 3222 14720
rect 3158 14660 3162 14716
rect 3162 14660 3218 14716
rect 3218 14660 3222 14716
rect 3158 14656 3222 14660
rect 6851 14716 6915 14720
rect 6851 14660 6855 14716
rect 6855 14660 6911 14716
rect 6911 14660 6915 14716
rect 6851 14656 6915 14660
rect 6931 14716 6995 14720
rect 6931 14660 6935 14716
rect 6935 14660 6991 14716
rect 6991 14660 6995 14716
rect 6931 14656 6995 14660
rect 7011 14716 7075 14720
rect 7011 14660 7015 14716
rect 7015 14660 7071 14716
rect 7071 14660 7075 14716
rect 7011 14656 7075 14660
rect 7091 14716 7155 14720
rect 7091 14660 7095 14716
rect 7095 14660 7151 14716
rect 7151 14660 7155 14716
rect 7091 14656 7155 14660
rect 10784 14716 10848 14720
rect 10784 14660 10788 14716
rect 10788 14660 10844 14716
rect 10844 14660 10848 14716
rect 10784 14656 10848 14660
rect 10864 14716 10928 14720
rect 10864 14660 10868 14716
rect 10868 14660 10924 14716
rect 10924 14660 10928 14716
rect 10864 14656 10928 14660
rect 10944 14716 11008 14720
rect 10944 14660 10948 14716
rect 10948 14660 11004 14716
rect 11004 14660 11008 14716
rect 10944 14656 11008 14660
rect 11024 14716 11088 14720
rect 11024 14660 11028 14716
rect 11028 14660 11084 14716
rect 11084 14660 11088 14716
rect 11024 14656 11088 14660
rect 14717 14716 14781 14720
rect 14717 14660 14721 14716
rect 14721 14660 14777 14716
rect 14777 14660 14781 14716
rect 14717 14656 14781 14660
rect 14797 14716 14861 14720
rect 14797 14660 14801 14716
rect 14801 14660 14857 14716
rect 14857 14660 14861 14716
rect 14797 14656 14861 14660
rect 14877 14716 14941 14720
rect 14877 14660 14881 14716
rect 14881 14660 14937 14716
rect 14937 14660 14941 14716
rect 14877 14656 14941 14660
rect 14957 14716 15021 14720
rect 14957 14660 14961 14716
rect 14961 14660 15017 14716
rect 15017 14660 15021 14716
rect 14957 14656 15021 14660
rect 4884 14172 4948 14176
rect 4884 14116 4888 14172
rect 4888 14116 4944 14172
rect 4944 14116 4948 14172
rect 4884 14112 4948 14116
rect 4964 14172 5028 14176
rect 4964 14116 4968 14172
rect 4968 14116 5024 14172
rect 5024 14116 5028 14172
rect 4964 14112 5028 14116
rect 5044 14172 5108 14176
rect 5044 14116 5048 14172
rect 5048 14116 5104 14172
rect 5104 14116 5108 14172
rect 5044 14112 5108 14116
rect 5124 14172 5188 14176
rect 5124 14116 5128 14172
rect 5128 14116 5184 14172
rect 5184 14116 5188 14172
rect 5124 14112 5188 14116
rect 8817 14172 8881 14176
rect 8817 14116 8821 14172
rect 8821 14116 8877 14172
rect 8877 14116 8881 14172
rect 8817 14112 8881 14116
rect 8897 14172 8961 14176
rect 8897 14116 8901 14172
rect 8901 14116 8957 14172
rect 8957 14116 8961 14172
rect 8897 14112 8961 14116
rect 8977 14172 9041 14176
rect 8977 14116 8981 14172
rect 8981 14116 9037 14172
rect 9037 14116 9041 14172
rect 8977 14112 9041 14116
rect 9057 14172 9121 14176
rect 9057 14116 9061 14172
rect 9061 14116 9117 14172
rect 9117 14116 9121 14172
rect 9057 14112 9121 14116
rect 12750 14172 12814 14176
rect 12750 14116 12754 14172
rect 12754 14116 12810 14172
rect 12810 14116 12814 14172
rect 12750 14112 12814 14116
rect 12830 14172 12894 14176
rect 12830 14116 12834 14172
rect 12834 14116 12890 14172
rect 12890 14116 12894 14172
rect 12830 14112 12894 14116
rect 12910 14172 12974 14176
rect 12910 14116 12914 14172
rect 12914 14116 12970 14172
rect 12970 14116 12974 14172
rect 12910 14112 12974 14116
rect 12990 14172 13054 14176
rect 12990 14116 12994 14172
rect 12994 14116 13050 14172
rect 13050 14116 13054 14172
rect 12990 14112 13054 14116
rect 16683 14172 16747 14176
rect 16683 14116 16687 14172
rect 16687 14116 16743 14172
rect 16743 14116 16747 14172
rect 16683 14112 16747 14116
rect 16763 14172 16827 14176
rect 16763 14116 16767 14172
rect 16767 14116 16823 14172
rect 16823 14116 16827 14172
rect 16763 14112 16827 14116
rect 16843 14172 16907 14176
rect 16843 14116 16847 14172
rect 16847 14116 16903 14172
rect 16903 14116 16907 14172
rect 16843 14112 16907 14116
rect 16923 14172 16987 14176
rect 16923 14116 16927 14172
rect 16927 14116 16983 14172
rect 16983 14116 16987 14172
rect 16923 14112 16987 14116
rect 2918 13628 2982 13632
rect 2918 13572 2922 13628
rect 2922 13572 2978 13628
rect 2978 13572 2982 13628
rect 2918 13568 2982 13572
rect 2998 13628 3062 13632
rect 2998 13572 3002 13628
rect 3002 13572 3058 13628
rect 3058 13572 3062 13628
rect 2998 13568 3062 13572
rect 3078 13628 3142 13632
rect 3078 13572 3082 13628
rect 3082 13572 3138 13628
rect 3138 13572 3142 13628
rect 3078 13568 3142 13572
rect 3158 13628 3222 13632
rect 3158 13572 3162 13628
rect 3162 13572 3218 13628
rect 3218 13572 3222 13628
rect 3158 13568 3222 13572
rect 6851 13628 6915 13632
rect 6851 13572 6855 13628
rect 6855 13572 6911 13628
rect 6911 13572 6915 13628
rect 6851 13568 6915 13572
rect 6931 13628 6995 13632
rect 6931 13572 6935 13628
rect 6935 13572 6991 13628
rect 6991 13572 6995 13628
rect 6931 13568 6995 13572
rect 7011 13628 7075 13632
rect 7011 13572 7015 13628
rect 7015 13572 7071 13628
rect 7071 13572 7075 13628
rect 7011 13568 7075 13572
rect 7091 13628 7155 13632
rect 7091 13572 7095 13628
rect 7095 13572 7151 13628
rect 7151 13572 7155 13628
rect 7091 13568 7155 13572
rect 10784 13628 10848 13632
rect 10784 13572 10788 13628
rect 10788 13572 10844 13628
rect 10844 13572 10848 13628
rect 10784 13568 10848 13572
rect 10864 13628 10928 13632
rect 10864 13572 10868 13628
rect 10868 13572 10924 13628
rect 10924 13572 10928 13628
rect 10864 13568 10928 13572
rect 10944 13628 11008 13632
rect 10944 13572 10948 13628
rect 10948 13572 11004 13628
rect 11004 13572 11008 13628
rect 10944 13568 11008 13572
rect 11024 13628 11088 13632
rect 11024 13572 11028 13628
rect 11028 13572 11084 13628
rect 11084 13572 11088 13628
rect 11024 13568 11088 13572
rect 14717 13628 14781 13632
rect 14717 13572 14721 13628
rect 14721 13572 14777 13628
rect 14777 13572 14781 13628
rect 14717 13568 14781 13572
rect 14797 13628 14861 13632
rect 14797 13572 14801 13628
rect 14801 13572 14857 13628
rect 14857 13572 14861 13628
rect 14797 13568 14861 13572
rect 14877 13628 14941 13632
rect 14877 13572 14881 13628
rect 14881 13572 14937 13628
rect 14937 13572 14941 13628
rect 14877 13568 14941 13572
rect 14957 13628 15021 13632
rect 14957 13572 14961 13628
rect 14961 13572 15017 13628
rect 15017 13572 15021 13628
rect 14957 13568 15021 13572
rect 4884 13084 4948 13088
rect 4884 13028 4888 13084
rect 4888 13028 4944 13084
rect 4944 13028 4948 13084
rect 4884 13024 4948 13028
rect 4964 13084 5028 13088
rect 4964 13028 4968 13084
rect 4968 13028 5024 13084
rect 5024 13028 5028 13084
rect 4964 13024 5028 13028
rect 5044 13084 5108 13088
rect 5044 13028 5048 13084
rect 5048 13028 5104 13084
rect 5104 13028 5108 13084
rect 5044 13024 5108 13028
rect 5124 13084 5188 13088
rect 5124 13028 5128 13084
rect 5128 13028 5184 13084
rect 5184 13028 5188 13084
rect 5124 13024 5188 13028
rect 8817 13084 8881 13088
rect 8817 13028 8821 13084
rect 8821 13028 8877 13084
rect 8877 13028 8881 13084
rect 8817 13024 8881 13028
rect 8897 13084 8961 13088
rect 8897 13028 8901 13084
rect 8901 13028 8957 13084
rect 8957 13028 8961 13084
rect 8897 13024 8961 13028
rect 8977 13084 9041 13088
rect 8977 13028 8981 13084
rect 8981 13028 9037 13084
rect 9037 13028 9041 13084
rect 8977 13024 9041 13028
rect 9057 13084 9121 13088
rect 9057 13028 9061 13084
rect 9061 13028 9117 13084
rect 9117 13028 9121 13084
rect 9057 13024 9121 13028
rect 12750 13084 12814 13088
rect 12750 13028 12754 13084
rect 12754 13028 12810 13084
rect 12810 13028 12814 13084
rect 12750 13024 12814 13028
rect 12830 13084 12894 13088
rect 12830 13028 12834 13084
rect 12834 13028 12890 13084
rect 12890 13028 12894 13084
rect 12830 13024 12894 13028
rect 12910 13084 12974 13088
rect 12910 13028 12914 13084
rect 12914 13028 12970 13084
rect 12970 13028 12974 13084
rect 12910 13024 12974 13028
rect 12990 13084 13054 13088
rect 12990 13028 12994 13084
rect 12994 13028 13050 13084
rect 13050 13028 13054 13084
rect 12990 13024 13054 13028
rect 16683 13084 16747 13088
rect 16683 13028 16687 13084
rect 16687 13028 16743 13084
rect 16743 13028 16747 13084
rect 16683 13024 16747 13028
rect 16763 13084 16827 13088
rect 16763 13028 16767 13084
rect 16767 13028 16823 13084
rect 16823 13028 16827 13084
rect 16763 13024 16827 13028
rect 16843 13084 16907 13088
rect 16843 13028 16847 13084
rect 16847 13028 16903 13084
rect 16903 13028 16907 13084
rect 16843 13024 16907 13028
rect 16923 13084 16987 13088
rect 16923 13028 16927 13084
rect 16927 13028 16983 13084
rect 16983 13028 16987 13084
rect 16923 13024 16987 13028
rect 2918 12540 2982 12544
rect 2918 12484 2922 12540
rect 2922 12484 2978 12540
rect 2978 12484 2982 12540
rect 2918 12480 2982 12484
rect 2998 12540 3062 12544
rect 2998 12484 3002 12540
rect 3002 12484 3058 12540
rect 3058 12484 3062 12540
rect 2998 12480 3062 12484
rect 3078 12540 3142 12544
rect 3078 12484 3082 12540
rect 3082 12484 3138 12540
rect 3138 12484 3142 12540
rect 3078 12480 3142 12484
rect 3158 12540 3222 12544
rect 3158 12484 3162 12540
rect 3162 12484 3218 12540
rect 3218 12484 3222 12540
rect 3158 12480 3222 12484
rect 6851 12540 6915 12544
rect 6851 12484 6855 12540
rect 6855 12484 6911 12540
rect 6911 12484 6915 12540
rect 6851 12480 6915 12484
rect 6931 12540 6995 12544
rect 6931 12484 6935 12540
rect 6935 12484 6991 12540
rect 6991 12484 6995 12540
rect 6931 12480 6995 12484
rect 7011 12540 7075 12544
rect 7011 12484 7015 12540
rect 7015 12484 7071 12540
rect 7071 12484 7075 12540
rect 7011 12480 7075 12484
rect 7091 12540 7155 12544
rect 7091 12484 7095 12540
rect 7095 12484 7151 12540
rect 7151 12484 7155 12540
rect 7091 12480 7155 12484
rect 10784 12540 10848 12544
rect 10784 12484 10788 12540
rect 10788 12484 10844 12540
rect 10844 12484 10848 12540
rect 10784 12480 10848 12484
rect 10864 12540 10928 12544
rect 10864 12484 10868 12540
rect 10868 12484 10924 12540
rect 10924 12484 10928 12540
rect 10864 12480 10928 12484
rect 10944 12540 11008 12544
rect 10944 12484 10948 12540
rect 10948 12484 11004 12540
rect 11004 12484 11008 12540
rect 10944 12480 11008 12484
rect 11024 12540 11088 12544
rect 11024 12484 11028 12540
rect 11028 12484 11084 12540
rect 11084 12484 11088 12540
rect 11024 12480 11088 12484
rect 14717 12540 14781 12544
rect 14717 12484 14721 12540
rect 14721 12484 14777 12540
rect 14777 12484 14781 12540
rect 14717 12480 14781 12484
rect 14797 12540 14861 12544
rect 14797 12484 14801 12540
rect 14801 12484 14857 12540
rect 14857 12484 14861 12540
rect 14797 12480 14861 12484
rect 14877 12540 14941 12544
rect 14877 12484 14881 12540
rect 14881 12484 14937 12540
rect 14937 12484 14941 12540
rect 14877 12480 14941 12484
rect 14957 12540 15021 12544
rect 14957 12484 14961 12540
rect 14961 12484 15017 12540
rect 15017 12484 15021 12540
rect 14957 12480 15021 12484
rect 4884 11996 4948 12000
rect 4884 11940 4888 11996
rect 4888 11940 4944 11996
rect 4944 11940 4948 11996
rect 4884 11936 4948 11940
rect 4964 11996 5028 12000
rect 4964 11940 4968 11996
rect 4968 11940 5024 11996
rect 5024 11940 5028 11996
rect 4964 11936 5028 11940
rect 5044 11996 5108 12000
rect 5044 11940 5048 11996
rect 5048 11940 5104 11996
rect 5104 11940 5108 11996
rect 5044 11936 5108 11940
rect 5124 11996 5188 12000
rect 5124 11940 5128 11996
rect 5128 11940 5184 11996
rect 5184 11940 5188 11996
rect 5124 11936 5188 11940
rect 8817 11996 8881 12000
rect 8817 11940 8821 11996
rect 8821 11940 8877 11996
rect 8877 11940 8881 11996
rect 8817 11936 8881 11940
rect 8897 11996 8961 12000
rect 8897 11940 8901 11996
rect 8901 11940 8957 11996
rect 8957 11940 8961 11996
rect 8897 11936 8961 11940
rect 8977 11996 9041 12000
rect 8977 11940 8981 11996
rect 8981 11940 9037 11996
rect 9037 11940 9041 11996
rect 8977 11936 9041 11940
rect 9057 11996 9121 12000
rect 9057 11940 9061 11996
rect 9061 11940 9117 11996
rect 9117 11940 9121 11996
rect 9057 11936 9121 11940
rect 12750 11996 12814 12000
rect 12750 11940 12754 11996
rect 12754 11940 12810 11996
rect 12810 11940 12814 11996
rect 12750 11936 12814 11940
rect 12830 11996 12894 12000
rect 12830 11940 12834 11996
rect 12834 11940 12890 11996
rect 12890 11940 12894 11996
rect 12830 11936 12894 11940
rect 12910 11996 12974 12000
rect 12910 11940 12914 11996
rect 12914 11940 12970 11996
rect 12970 11940 12974 11996
rect 12910 11936 12974 11940
rect 12990 11996 13054 12000
rect 12990 11940 12994 11996
rect 12994 11940 13050 11996
rect 13050 11940 13054 11996
rect 12990 11936 13054 11940
rect 16683 11996 16747 12000
rect 16683 11940 16687 11996
rect 16687 11940 16743 11996
rect 16743 11940 16747 11996
rect 16683 11936 16747 11940
rect 16763 11996 16827 12000
rect 16763 11940 16767 11996
rect 16767 11940 16823 11996
rect 16823 11940 16827 11996
rect 16763 11936 16827 11940
rect 16843 11996 16907 12000
rect 16843 11940 16847 11996
rect 16847 11940 16903 11996
rect 16903 11940 16907 11996
rect 16843 11936 16907 11940
rect 16923 11996 16987 12000
rect 16923 11940 16927 11996
rect 16927 11940 16983 11996
rect 16983 11940 16987 11996
rect 16923 11936 16987 11940
rect 2918 11452 2982 11456
rect 2918 11396 2922 11452
rect 2922 11396 2978 11452
rect 2978 11396 2982 11452
rect 2918 11392 2982 11396
rect 2998 11452 3062 11456
rect 2998 11396 3002 11452
rect 3002 11396 3058 11452
rect 3058 11396 3062 11452
rect 2998 11392 3062 11396
rect 3078 11452 3142 11456
rect 3078 11396 3082 11452
rect 3082 11396 3138 11452
rect 3138 11396 3142 11452
rect 3078 11392 3142 11396
rect 3158 11452 3222 11456
rect 3158 11396 3162 11452
rect 3162 11396 3218 11452
rect 3218 11396 3222 11452
rect 3158 11392 3222 11396
rect 6851 11452 6915 11456
rect 6851 11396 6855 11452
rect 6855 11396 6911 11452
rect 6911 11396 6915 11452
rect 6851 11392 6915 11396
rect 6931 11452 6995 11456
rect 6931 11396 6935 11452
rect 6935 11396 6991 11452
rect 6991 11396 6995 11452
rect 6931 11392 6995 11396
rect 7011 11452 7075 11456
rect 7011 11396 7015 11452
rect 7015 11396 7071 11452
rect 7071 11396 7075 11452
rect 7011 11392 7075 11396
rect 7091 11452 7155 11456
rect 7091 11396 7095 11452
rect 7095 11396 7151 11452
rect 7151 11396 7155 11452
rect 7091 11392 7155 11396
rect 10784 11452 10848 11456
rect 10784 11396 10788 11452
rect 10788 11396 10844 11452
rect 10844 11396 10848 11452
rect 10784 11392 10848 11396
rect 10864 11452 10928 11456
rect 10864 11396 10868 11452
rect 10868 11396 10924 11452
rect 10924 11396 10928 11452
rect 10864 11392 10928 11396
rect 10944 11452 11008 11456
rect 10944 11396 10948 11452
rect 10948 11396 11004 11452
rect 11004 11396 11008 11452
rect 10944 11392 11008 11396
rect 11024 11452 11088 11456
rect 11024 11396 11028 11452
rect 11028 11396 11084 11452
rect 11084 11396 11088 11452
rect 11024 11392 11088 11396
rect 14717 11452 14781 11456
rect 14717 11396 14721 11452
rect 14721 11396 14777 11452
rect 14777 11396 14781 11452
rect 14717 11392 14781 11396
rect 14797 11452 14861 11456
rect 14797 11396 14801 11452
rect 14801 11396 14857 11452
rect 14857 11396 14861 11452
rect 14797 11392 14861 11396
rect 14877 11452 14941 11456
rect 14877 11396 14881 11452
rect 14881 11396 14937 11452
rect 14937 11396 14941 11452
rect 14877 11392 14941 11396
rect 14957 11452 15021 11456
rect 14957 11396 14961 11452
rect 14961 11396 15017 11452
rect 15017 11396 15021 11452
rect 14957 11392 15021 11396
rect 4884 10908 4948 10912
rect 4884 10852 4888 10908
rect 4888 10852 4944 10908
rect 4944 10852 4948 10908
rect 4884 10848 4948 10852
rect 4964 10908 5028 10912
rect 4964 10852 4968 10908
rect 4968 10852 5024 10908
rect 5024 10852 5028 10908
rect 4964 10848 5028 10852
rect 5044 10908 5108 10912
rect 5044 10852 5048 10908
rect 5048 10852 5104 10908
rect 5104 10852 5108 10908
rect 5044 10848 5108 10852
rect 5124 10908 5188 10912
rect 5124 10852 5128 10908
rect 5128 10852 5184 10908
rect 5184 10852 5188 10908
rect 5124 10848 5188 10852
rect 8817 10908 8881 10912
rect 8817 10852 8821 10908
rect 8821 10852 8877 10908
rect 8877 10852 8881 10908
rect 8817 10848 8881 10852
rect 8897 10908 8961 10912
rect 8897 10852 8901 10908
rect 8901 10852 8957 10908
rect 8957 10852 8961 10908
rect 8897 10848 8961 10852
rect 8977 10908 9041 10912
rect 8977 10852 8981 10908
rect 8981 10852 9037 10908
rect 9037 10852 9041 10908
rect 8977 10848 9041 10852
rect 9057 10908 9121 10912
rect 9057 10852 9061 10908
rect 9061 10852 9117 10908
rect 9117 10852 9121 10908
rect 9057 10848 9121 10852
rect 12750 10908 12814 10912
rect 12750 10852 12754 10908
rect 12754 10852 12810 10908
rect 12810 10852 12814 10908
rect 12750 10848 12814 10852
rect 12830 10908 12894 10912
rect 12830 10852 12834 10908
rect 12834 10852 12890 10908
rect 12890 10852 12894 10908
rect 12830 10848 12894 10852
rect 12910 10908 12974 10912
rect 12910 10852 12914 10908
rect 12914 10852 12970 10908
rect 12970 10852 12974 10908
rect 12910 10848 12974 10852
rect 12990 10908 13054 10912
rect 12990 10852 12994 10908
rect 12994 10852 13050 10908
rect 13050 10852 13054 10908
rect 12990 10848 13054 10852
rect 16683 10908 16747 10912
rect 16683 10852 16687 10908
rect 16687 10852 16743 10908
rect 16743 10852 16747 10908
rect 16683 10848 16747 10852
rect 16763 10908 16827 10912
rect 16763 10852 16767 10908
rect 16767 10852 16823 10908
rect 16823 10852 16827 10908
rect 16763 10848 16827 10852
rect 16843 10908 16907 10912
rect 16843 10852 16847 10908
rect 16847 10852 16903 10908
rect 16903 10852 16907 10908
rect 16843 10848 16907 10852
rect 16923 10908 16987 10912
rect 16923 10852 16927 10908
rect 16927 10852 16983 10908
rect 16983 10852 16987 10908
rect 16923 10848 16987 10852
rect 2918 10364 2982 10368
rect 2918 10308 2922 10364
rect 2922 10308 2978 10364
rect 2978 10308 2982 10364
rect 2918 10304 2982 10308
rect 2998 10364 3062 10368
rect 2998 10308 3002 10364
rect 3002 10308 3058 10364
rect 3058 10308 3062 10364
rect 2998 10304 3062 10308
rect 3078 10364 3142 10368
rect 3078 10308 3082 10364
rect 3082 10308 3138 10364
rect 3138 10308 3142 10364
rect 3078 10304 3142 10308
rect 3158 10364 3222 10368
rect 3158 10308 3162 10364
rect 3162 10308 3218 10364
rect 3218 10308 3222 10364
rect 3158 10304 3222 10308
rect 6851 10364 6915 10368
rect 6851 10308 6855 10364
rect 6855 10308 6911 10364
rect 6911 10308 6915 10364
rect 6851 10304 6915 10308
rect 6931 10364 6995 10368
rect 6931 10308 6935 10364
rect 6935 10308 6991 10364
rect 6991 10308 6995 10364
rect 6931 10304 6995 10308
rect 7011 10364 7075 10368
rect 7011 10308 7015 10364
rect 7015 10308 7071 10364
rect 7071 10308 7075 10364
rect 7011 10304 7075 10308
rect 7091 10364 7155 10368
rect 7091 10308 7095 10364
rect 7095 10308 7151 10364
rect 7151 10308 7155 10364
rect 7091 10304 7155 10308
rect 10784 10364 10848 10368
rect 10784 10308 10788 10364
rect 10788 10308 10844 10364
rect 10844 10308 10848 10364
rect 10784 10304 10848 10308
rect 10864 10364 10928 10368
rect 10864 10308 10868 10364
rect 10868 10308 10924 10364
rect 10924 10308 10928 10364
rect 10864 10304 10928 10308
rect 10944 10364 11008 10368
rect 10944 10308 10948 10364
rect 10948 10308 11004 10364
rect 11004 10308 11008 10364
rect 10944 10304 11008 10308
rect 11024 10364 11088 10368
rect 11024 10308 11028 10364
rect 11028 10308 11084 10364
rect 11084 10308 11088 10364
rect 11024 10304 11088 10308
rect 14717 10364 14781 10368
rect 14717 10308 14721 10364
rect 14721 10308 14777 10364
rect 14777 10308 14781 10364
rect 14717 10304 14781 10308
rect 14797 10364 14861 10368
rect 14797 10308 14801 10364
rect 14801 10308 14857 10364
rect 14857 10308 14861 10364
rect 14797 10304 14861 10308
rect 14877 10364 14941 10368
rect 14877 10308 14881 10364
rect 14881 10308 14937 10364
rect 14937 10308 14941 10364
rect 14877 10304 14941 10308
rect 14957 10364 15021 10368
rect 14957 10308 14961 10364
rect 14961 10308 15017 10364
rect 15017 10308 15021 10364
rect 14957 10304 15021 10308
rect 4884 9820 4948 9824
rect 4884 9764 4888 9820
rect 4888 9764 4944 9820
rect 4944 9764 4948 9820
rect 4884 9760 4948 9764
rect 4964 9820 5028 9824
rect 4964 9764 4968 9820
rect 4968 9764 5024 9820
rect 5024 9764 5028 9820
rect 4964 9760 5028 9764
rect 5044 9820 5108 9824
rect 5044 9764 5048 9820
rect 5048 9764 5104 9820
rect 5104 9764 5108 9820
rect 5044 9760 5108 9764
rect 5124 9820 5188 9824
rect 5124 9764 5128 9820
rect 5128 9764 5184 9820
rect 5184 9764 5188 9820
rect 5124 9760 5188 9764
rect 8817 9820 8881 9824
rect 8817 9764 8821 9820
rect 8821 9764 8877 9820
rect 8877 9764 8881 9820
rect 8817 9760 8881 9764
rect 8897 9820 8961 9824
rect 8897 9764 8901 9820
rect 8901 9764 8957 9820
rect 8957 9764 8961 9820
rect 8897 9760 8961 9764
rect 8977 9820 9041 9824
rect 8977 9764 8981 9820
rect 8981 9764 9037 9820
rect 9037 9764 9041 9820
rect 8977 9760 9041 9764
rect 9057 9820 9121 9824
rect 9057 9764 9061 9820
rect 9061 9764 9117 9820
rect 9117 9764 9121 9820
rect 9057 9760 9121 9764
rect 12750 9820 12814 9824
rect 12750 9764 12754 9820
rect 12754 9764 12810 9820
rect 12810 9764 12814 9820
rect 12750 9760 12814 9764
rect 12830 9820 12894 9824
rect 12830 9764 12834 9820
rect 12834 9764 12890 9820
rect 12890 9764 12894 9820
rect 12830 9760 12894 9764
rect 12910 9820 12974 9824
rect 12910 9764 12914 9820
rect 12914 9764 12970 9820
rect 12970 9764 12974 9820
rect 12910 9760 12974 9764
rect 12990 9820 13054 9824
rect 12990 9764 12994 9820
rect 12994 9764 13050 9820
rect 13050 9764 13054 9820
rect 12990 9760 13054 9764
rect 16683 9820 16747 9824
rect 16683 9764 16687 9820
rect 16687 9764 16743 9820
rect 16743 9764 16747 9820
rect 16683 9760 16747 9764
rect 16763 9820 16827 9824
rect 16763 9764 16767 9820
rect 16767 9764 16823 9820
rect 16823 9764 16827 9820
rect 16763 9760 16827 9764
rect 16843 9820 16907 9824
rect 16843 9764 16847 9820
rect 16847 9764 16903 9820
rect 16903 9764 16907 9820
rect 16843 9760 16907 9764
rect 16923 9820 16987 9824
rect 16923 9764 16927 9820
rect 16927 9764 16983 9820
rect 16983 9764 16987 9820
rect 16923 9760 16987 9764
rect 2918 9276 2982 9280
rect 2918 9220 2922 9276
rect 2922 9220 2978 9276
rect 2978 9220 2982 9276
rect 2918 9216 2982 9220
rect 2998 9276 3062 9280
rect 2998 9220 3002 9276
rect 3002 9220 3058 9276
rect 3058 9220 3062 9276
rect 2998 9216 3062 9220
rect 3078 9276 3142 9280
rect 3078 9220 3082 9276
rect 3082 9220 3138 9276
rect 3138 9220 3142 9276
rect 3078 9216 3142 9220
rect 3158 9276 3222 9280
rect 3158 9220 3162 9276
rect 3162 9220 3218 9276
rect 3218 9220 3222 9276
rect 3158 9216 3222 9220
rect 6851 9276 6915 9280
rect 6851 9220 6855 9276
rect 6855 9220 6911 9276
rect 6911 9220 6915 9276
rect 6851 9216 6915 9220
rect 6931 9276 6995 9280
rect 6931 9220 6935 9276
rect 6935 9220 6991 9276
rect 6991 9220 6995 9276
rect 6931 9216 6995 9220
rect 7011 9276 7075 9280
rect 7011 9220 7015 9276
rect 7015 9220 7071 9276
rect 7071 9220 7075 9276
rect 7011 9216 7075 9220
rect 7091 9276 7155 9280
rect 7091 9220 7095 9276
rect 7095 9220 7151 9276
rect 7151 9220 7155 9276
rect 7091 9216 7155 9220
rect 10784 9276 10848 9280
rect 10784 9220 10788 9276
rect 10788 9220 10844 9276
rect 10844 9220 10848 9276
rect 10784 9216 10848 9220
rect 10864 9276 10928 9280
rect 10864 9220 10868 9276
rect 10868 9220 10924 9276
rect 10924 9220 10928 9276
rect 10864 9216 10928 9220
rect 10944 9276 11008 9280
rect 10944 9220 10948 9276
rect 10948 9220 11004 9276
rect 11004 9220 11008 9276
rect 10944 9216 11008 9220
rect 11024 9276 11088 9280
rect 11024 9220 11028 9276
rect 11028 9220 11084 9276
rect 11084 9220 11088 9276
rect 11024 9216 11088 9220
rect 14717 9276 14781 9280
rect 14717 9220 14721 9276
rect 14721 9220 14777 9276
rect 14777 9220 14781 9276
rect 14717 9216 14781 9220
rect 14797 9276 14861 9280
rect 14797 9220 14801 9276
rect 14801 9220 14857 9276
rect 14857 9220 14861 9276
rect 14797 9216 14861 9220
rect 14877 9276 14941 9280
rect 14877 9220 14881 9276
rect 14881 9220 14937 9276
rect 14937 9220 14941 9276
rect 14877 9216 14941 9220
rect 14957 9276 15021 9280
rect 14957 9220 14961 9276
rect 14961 9220 15017 9276
rect 15017 9220 15021 9276
rect 14957 9216 15021 9220
rect 4884 8732 4948 8736
rect 4884 8676 4888 8732
rect 4888 8676 4944 8732
rect 4944 8676 4948 8732
rect 4884 8672 4948 8676
rect 4964 8732 5028 8736
rect 4964 8676 4968 8732
rect 4968 8676 5024 8732
rect 5024 8676 5028 8732
rect 4964 8672 5028 8676
rect 5044 8732 5108 8736
rect 5044 8676 5048 8732
rect 5048 8676 5104 8732
rect 5104 8676 5108 8732
rect 5044 8672 5108 8676
rect 5124 8732 5188 8736
rect 5124 8676 5128 8732
rect 5128 8676 5184 8732
rect 5184 8676 5188 8732
rect 5124 8672 5188 8676
rect 8817 8732 8881 8736
rect 8817 8676 8821 8732
rect 8821 8676 8877 8732
rect 8877 8676 8881 8732
rect 8817 8672 8881 8676
rect 8897 8732 8961 8736
rect 8897 8676 8901 8732
rect 8901 8676 8957 8732
rect 8957 8676 8961 8732
rect 8897 8672 8961 8676
rect 8977 8732 9041 8736
rect 8977 8676 8981 8732
rect 8981 8676 9037 8732
rect 9037 8676 9041 8732
rect 8977 8672 9041 8676
rect 9057 8732 9121 8736
rect 9057 8676 9061 8732
rect 9061 8676 9117 8732
rect 9117 8676 9121 8732
rect 9057 8672 9121 8676
rect 12750 8732 12814 8736
rect 12750 8676 12754 8732
rect 12754 8676 12810 8732
rect 12810 8676 12814 8732
rect 12750 8672 12814 8676
rect 12830 8732 12894 8736
rect 12830 8676 12834 8732
rect 12834 8676 12890 8732
rect 12890 8676 12894 8732
rect 12830 8672 12894 8676
rect 12910 8732 12974 8736
rect 12910 8676 12914 8732
rect 12914 8676 12970 8732
rect 12970 8676 12974 8732
rect 12910 8672 12974 8676
rect 12990 8732 13054 8736
rect 12990 8676 12994 8732
rect 12994 8676 13050 8732
rect 13050 8676 13054 8732
rect 12990 8672 13054 8676
rect 16683 8732 16747 8736
rect 16683 8676 16687 8732
rect 16687 8676 16743 8732
rect 16743 8676 16747 8732
rect 16683 8672 16747 8676
rect 16763 8732 16827 8736
rect 16763 8676 16767 8732
rect 16767 8676 16823 8732
rect 16823 8676 16827 8732
rect 16763 8672 16827 8676
rect 16843 8732 16907 8736
rect 16843 8676 16847 8732
rect 16847 8676 16903 8732
rect 16903 8676 16907 8732
rect 16843 8672 16907 8676
rect 16923 8732 16987 8736
rect 16923 8676 16927 8732
rect 16927 8676 16983 8732
rect 16983 8676 16987 8732
rect 16923 8672 16987 8676
rect 2918 8188 2982 8192
rect 2918 8132 2922 8188
rect 2922 8132 2978 8188
rect 2978 8132 2982 8188
rect 2918 8128 2982 8132
rect 2998 8188 3062 8192
rect 2998 8132 3002 8188
rect 3002 8132 3058 8188
rect 3058 8132 3062 8188
rect 2998 8128 3062 8132
rect 3078 8188 3142 8192
rect 3078 8132 3082 8188
rect 3082 8132 3138 8188
rect 3138 8132 3142 8188
rect 3078 8128 3142 8132
rect 3158 8188 3222 8192
rect 3158 8132 3162 8188
rect 3162 8132 3218 8188
rect 3218 8132 3222 8188
rect 3158 8128 3222 8132
rect 6851 8188 6915 8192
rect 6851 8132 6855 8188
rect 6855 8132 6911 8188
rect 6911 8132 6915 8188
rect 6851 8128 6915 8132
rect 6931 8188 6995 8192
rect 6931 8132 6935 8188
rect 6935 8132 6991 8188
rect 6991 8132 6995 8188
rect 6931 8128 6995 8132
rect 7011 8188 7075 8192
rect 7011 8132 7015 8188
rect 7015 8132 7071 8188
rect 7071 8132 7075 8188
rect 7011 8128 7075 8132
rect 7091 8188 7155 8192
rect 7091 8132 7095 8188
rect 7095 8132 7151 8188
rect 7151 8132 7155 8188
rect 7091 8128 7155 8132
rect 10784 8188 10848 8192
rect 10784 8132 10788 8188
rect 10788 8132 10844 8188
rect 10844 8132 10848 8188
rect 10784 8128 10848 8132
rect 10864 8188 10928 8192
rect 10864 8132 10868 8188
rect 10868 8132 10924 8188
rect 10924 8132 10928 8188
rect 10864 8128 10928 8132
rect 10944 8188 11008 8192
rect 10944 8132 10948 8188
rect 10948 8132 11004 8188
rect 11004 8132 11008 8188
rect 10944 8128 11008 8132
rect 11024 8188 11088 8192
rect 11024 8132 11028 8188
rect 11028 8132 11084 8188
rect 11084 8132 11088 8188
rect 11024 8128 11088 8132
rect 14717 8188 14781 8192
rect 14717 8132 14721 8188
rect 14721 8132 14777 8188
rect 14777 8132 14781 8188
rect 14717 8128 14781 8132
rect 14797 8188 14861 8192
rect 14797 8132 14801 8188
rect 14801 8132 14857 8188
rect 14857 8132 14861 8188
rect 14797 8128 14861 8132
rect 14877 8188 14941 8192
rect 14877 8132 14881 8188
rect 14881 8132 14937 8188
rect 14937 8132 14941 8188
rect 14877 8128 14941 8132
rect 14957 8188 15021 8192
rect 14957 8132 14961 8188
rect 14961 8132 15017 8188
rect 15017 8132 15021 8188
rect 14957 8128 15021 8132
rect 4884 7644 4948 7648
rect 4884 7588 4888 7644
rect 4888 7588 4944 7644
rect 4944 7588 4948 7644
rect 4884 7584 4948 7588
rect 4964 7644 5028 7648
rect 4964 7588 4968 7644
rect 4968 7588 5024 7644
rect 5024 7588 5028 7644
rect 4964 7584 5028 7588
rect 5044 7644 5108 7648
rect 5044 7588 5048 7644
rect 5048 7588 5104 7644
rect 5104 7588 5108 7644
rect 5044 7584 5108 7588
rect 5124 7644 5188 7648
rect 5124 7588 5128 7644
rect 5128 7588 5184 7644
rect 5184 7588 5188 7644
rect 5124 7584 5188 7588
rect 8817 7644 8881 7648
rect 8817 7588 8821 7644
rect 8821 7588 8877 7644
rect 8877 7588 8881 7644
rect 8817 7584 8881 7588
rect 8897 7644 8961 7648
rect 8897 7588 8901 7644
rect 8901 7588 8957 7644
rect 8957 7588 8961 7644
rect 8897 7584 8961 7588
rect 8977 7644 9041 7648
rect 8977 7588 8981 7644
rect 8981 7588 9037 7644
rect 9037 7588 9041 7644
rect 8977 7584 9041 7588
rect 9057 7644 9121 7648
rect 9057 7588 9061 7644
rect 9061 7588 9117 7644
rect 9117 7588 9121 7644
rect 9057 7584 9121 7588
rect 12750 7644 12814 7648
rect 12750 7588 12754 7644
rect 12754 7588 12810 7644
rect 12810 7588 12814 7644
rect 12750 7584 12814 7588
rect 12830 7644 12894 7648
rect 12830 7588 12834 7644
rect 12834 7588 12890 7644
rect 12890 7588 12894 7644
rect 12830 7584 12894 7588
rect 12910 7644 12974 7648
rect 12910 7588 12914 7644
rect 12914 7588 12970 7644
rect 12970 7588 12974 7644
rect 12910 7584 12974 7588
rect 12990 7644 13054 7648
rect 12990 7588 12994 7644
rect 12994 7588 13050 7644
rect 13050 7588 13054 7644
rect 12990 7584 13054 7588
rect 16683 7644 16747 7648
rect 16683 7588 16687 7644
rect 16687 7588 16743 7644
rect 16743 7588 16747 7644
rect 16683 7584 16747 7588
rect 16763 7644 16827 7648
rect 16763 7588 16767 7644
rect 16767 7588 16823 7644
rect 16823 7588 16827 7644
rect 16763 7584 16827 7588
rect 16843 7644 16907 7648
rect 16843 7588 16847 7644
rect 16847 7588 16903 7644
rect 16903 7588 16907 7644
rect 16843 7584 16907 7588
rect 16923 7644 16987 7648
rect 16923 7588 16927 7644
rect 16927 7588 16983 7644
rect 16983 7588 16987 7644
rect 16923 7584 16987 7588
rect 2918 7100 2982 7104
rect 2918 7044 2922 7100
rect 2922 7044 2978 7100
rect 2978 7044 2982 7100
rect 2918 7040 2982 7044
rect 2998 7100 3062 7104
rect 2998 7044 3002 7100
rect 3002 7044 3058 7100
rect 3058 7044 3062 7100
rect 2998 7040 3062 7044
rect 3078 7100 3142 7104
rect 3078 7044 3082 7100
rect 3082 7044 3138 7100
rect 3138 7044 3142 7100
rect 3078 7040 3142 7044
rect 3158 7100 3222 7104
rect 3158 7044 3162 7100
rect 3162 7044 3218 7100
rect 3218 7044 3222 7100
rect 3158 7040 3222 7044
rect 6851 7100 6915 7104
rect 6851 7044 6855 7100
rect 6855 7044 6911 7100
rect 6911 7044 6915 7100
rect 6851 7040 6915 7044
rect 6931 7100 6995 7104
rect 6931 7044 6935 7100
rect 6935 7044 6991 7100
rect 6991 7044 6995 7100
rect 6931 7040 6995 7044
rect 7011 7100 7075 7104
rect 7011 7044 7015 7100
rect 7015 7044 7071 7100
rect 7071 7044 7075 7100
rect 7011 7040 7075 7044
rect 7091 7100 7155 7104
rect 7091 7044 7095 7100
rect 7095 7044 7151 7100
rect 7151 7044 7155 7100
rect 7091 7040 7155 7044
rect 10784 7100 10848 7104
rect 10784 7044 10788 7100
rect 10788 7044 10844 7100
rect 10844 7044 10848 7100
rect 10784 7040 10848 7044
rect 10864 7100 10928 7104
rect 10864 7044 10868 7100
rect 10868 7044 10924 7100
rect 10924 7044 10928 7100
rect 10864 7040 10928 7044
rect 10944 7100 11008 7104
rect 10944 7044 10948 7100
rect 10948 7044 11004 7100
rect 11004 7044 11008 7100
rect 10944 7040 11008 7044
rect 11024 7100 11088 7104
rect 11024 7044 11028 7100
rect 11028 7044 11084 7100
rect 11084 7044 11088 7100
rect 11024 7040 11088 7044
rect 14717 7100 14781 7104
rect 14717 7044 14721 7100
rect 14721 7044 14777 7100
rect 14777 7044 14781 7100
rect 14717 7040 14781 7044
rect 14797 7100 14861 7104
rect 14797 7044 14801 7100
rect 14801 7044 14857 7100
rect 14857 7044 14861 7100
rect 14797 7040 14861 7044
rect 14877 7100 14941 7104
rect 14877 7044 14881 7100
rect 14881 7044 14937 7100
rect 14937 7044 14941 7100
rect 14877 7040 14941 7044
rect 14957 7100 15021 7104
rect 14957 7044 14961 7100
rect 14961 7044 15017 7100
rect 15017 7044 15021 7100
rect 14957 7040 15021 7044
rect 4884 6556 4948 6560
rect 4884 6500 4888 6556
rect 4888 6500 4944 6556
rect 4944 6500 4948 6556
rect 4884 6496 4948 6500
rect 4964 6556 5028 6560
rect 4964 6500 4968 6556
rect 4968 6500 5024 6556
rect 5024 6500 5028 6556
rect 4964 6496 5028 6500
rect 5044 6556 5108 6560
rect 5044 6500 5048 6556
rect 5048 6500 5104 6556
rect 5104 6500 5108 6556
rect 5044 6496 5108 6500
rect 5124 6556 5188 6560
rect 5124 6500 5128 6556
rect 5128 6500 5184 6556
rect 5184 6500 5188 6556
rect 5124 6496 5188 6500
rect 8817 6556 8881 6560
rect 8817 6500 8821 6556
rect 8821 6500 8877 6556
rect 8877 6500 8881 6556
rect 8817 6496 8881 6500
rect 8897 6556 8961 6560
rect 8897 6500 8901 6556
rect 8901 6500 8957 6556
rect 8957 6500 8961 6556
rect 8897 6496 8961 6500
rect 8977 6556 9041 6560
rect 8977 6500 8981 6556
rect 8981 6500 9037 6556
rect 9037 6500 9041 6556
rect 8977 6496 9041 6500
rect 9057 6556 9121 6560
rect 9057 6500 9061 6556
rect 9061 6500 9117 6556
rect 9117 6500 9121 6556
rect 9057 6496 9121 6500
rect 12750 6556 12814 6560
rect 12750 6500 12754 6556
rect 12754 6500 12810 6556
rect 12810 6500 12814 6556
rect 12750 6496 12814 6500
rect 12830 6556 12894 6560
rect 12830 6500 12834 6556
rect 12834 6500 12890 6556
rect 12890 6500 12894 6556
rect 12830 6496 12894 6500
rect 12910 6556 12974 6560
rect 12910 6500 12914 6556
rect 12914 6500 12970 6556
rect 12970 6500 12974 6556
rect 12910 6496 12974 6500
rect 12990 6556 13054 6560
rect 12990 6500 12994 6556
rect 12994 6500 13050 6556
rect 13050 6500 13054 6556
rect 12990 6496 13054 6500
rect 16683 6556 16747 6560
rect 16683 6500 16687 6556
rect 16687 6500 16743 6556
rect 16743 6500 16747 6556
rect 16683 6496 16747 6500
rect 16763 6556 16827 6560
rect 16763 6500 16767 6556
rect 16767 6500 16823 6556
rect 16823 6500 16827 6556
rect 16763 6496 16827 6500
rect 16843 6556 16907 6560
rect 16843 6500 16847 6556
rect 16847 6500 16903 6556
rect 16903 6500 16907 6556
rect 16843 6496 16907 6500
rect 16923 6556 16987 6560
rect 16923 6500 16927 6556
rect 16927 6500 16983 6556
rect 16983 6500 16987 6556
rect 16923 6496 16987 6500
rect 2918 6012 2982 6016
rect 2918 5956 2922 6012
rect 2922 5956 2978 6012
rect 2978 5956 2982 6012
rect 2918 5952 2982 5956
rect 2998 6012 3062 6016
rect 2998 5956 3002 6012
rect 3002 5956 3058 6012
rect 3058 5956 3062 6012
rect 2998 5952 3062 5956
rect 3078 6012 3142 6016
rect 3078 5956 3082 6012
rect 3082 5956 3138 6012
rect 3138 5956 3142 6012
rect 3078 5952 3142 5956
rect 3158 6012 3222 6016
rect 3158 5956 3162 6012
rect 3162 5956 3218 6012
rect 3218 5956 3222 6012
rect 3158 5952 3222 5956
rect 6851 6012 6915 6016
rect 6851 5956 6855 6012
rect 6855 5956 6911 6012
rect 6911 5956 6915 6012
rect 6851 5952 6915 5956
rect 6931 6012 6995 6016
rect 6931 5956 6935 6012
rect 6935 5956 6991 6012
rect 6991 5956 6995 6012
rect 6931 5952 6995 5956
rect 7011 6012 7075 6016
rect 7011 5956 7015 6012
rect 7015 5956 7071 6012
rect 7071 5956 7075 6012
rect 7011 5952 7075 5956
rect 7091 6012 7155 6016
rect 7091 5956 7095 6012
rect 7095 5956 7151 6012
rect 7151 5956 7155 6012
rect 7091 5952 7155 5956
rect 10784 6012 10848 6016
rect 10784 5956 10788 6012
rect 10788 5956 10844 6012
rect 10844 5956 10848 6012
rect 10784 5952 10848 5956
rect 10864 6012 10928 6016
rect 10864 5956 10868 6012
rect 10868 5956 10924 6012
rect 10924 5956 10928 6012
rect 10864 5952 10928 5956
rect 10944 6012 11008 6016
rect 10944 5956 10948 6012
rect 10948 5956 11004 6012
rect 11004 5956 11008 6012
rect 10944 5952 11008 5956
rect 11024 6012 11088 6016
rect 11024 5956 11028 6012
rect 11028 5956 11084 6012
rect 11084 5956 11088 6012
rect 11024 5952 11088 5956
rect 14717 6012 14781 6016
rect 14717 5956 14721 6012
rect 14721 5956 14777 6012
rect 14777 5956 14781 6012
rect 14717 5952 14781 5956
rect 14797 6012 14861 6016
rect 14797 5956 14801 6012
rect 14801 5956 14857 6012
rect 14857 5956 14861 6012
rect 14797 5952 14861 5956
rect 14877 6012 14941 6016
rect 14877 5956 14881 6012
rect 14881 5956 14937 6012
rect 14937 5956 14941 6012
rect 14877 5952 14941 5956
rect 14957 6012 15021 6016
rect 14957 5956 14961 6012
rect 14961 5956 15017 6012
rect 15017 5956 15021 6012
rect 14957 5952 15021 5956
rect 4884 5468 4948 5472
rect 4884 5412 4888 5468
rect 4888 5412 4944 5468
rect 4944 5412 4948 5468
rect 4884 5408 4948 5412
rect 4964 5468 5028 5472
rect 4964 5412 4968 5468
rect 4968 5412 5024 5468
rect 5024 5412 5028 5468
rect 4964 5408 5028 5412
rect 5044 5468 5108 5472
rect 5044 5412 5048 5468
rect 5048 5412 5104 5468
rect 5104 5412 5108 5468
rect 5044 5408 5108 5412
rect 5124 5468 5188 5472
rect 5124 5412 5128 5468
rect 5128 5412 5184 5468
rect 5184 5412 5188 5468
rect 5124 5408 5188 5412
rect 8817 5468 8881 5472
rect 8817 5412 8821 5468
rect 8821 5412 8877 5468
rect 8877 5412 8881 5468
rect 8817 5408 8881 5412
rect 8897 5468 8961 5472
rect 8897 5412 8901 5468
rect 8901 5412 8957 5468
rect 8957 5412 8961 5468
rect 8897 5408 8961 5412
rect 8977 5468 9041 5472
rect 8977 5412 8981 5468
rect 8981 5412 9037 5468
rect 9037 5412 9041 5468
rect 8977 5408 9041 5412
rect 9057 5468 9121 5472
rect 9057 5412 9061 5468
rect 9061 5412 9117 5468
rect 9117 5412 9121 5468
rect 9057 5408 9121 5412
rect 12750 5468 12814 5472
rect 12750 5412 12754 5468
rect 12754 5412 12810 5468
rect 12810 5412 12814 5468
rect 12750 5408 12814 5412
rect 12830 5468 12894 5472
rect 12830 5412 12834 5468
rect 12834 5412 12890 5468
rect 12890 5412 12894 5468
rect 12830 5408 12894 5412
rect 12910 5468 12974 5472
rect 12910 5412 12914 5468
rect 12914 5412 12970 5468
rect 12970 5412 12974 5468
rect 12910 5408 12974 5412
rect 12990 5468 13054 5472
rect 12990 5412 12994 5468
rect 12994 5412 13050 5468
rect 13050 5412 13054 5468
rect 12990 5408 13054 5412
rect 16683 5468 16747 5472
rect 16683 5412 16687 5468
rect 16687 5412 16743 5468
rect 16743 5412 16747 5468
rect 16683 5408 16747 5412
rect 16763 5468 16827 5472
rect 16763 5412 16767 5468
rect 16767 5412 16823 5468
rect 16823 5412 16827 5468
rect 16763 5408 16827 5412
rect 16843 5468 16907 5472
rect 16843 5412 16847 5468
rect 16847 5412 16903 5468
rect 16903 5412 16907 5468
rect 16843 5408 16907 5412
rect 16923 5468 16987 5472
rect 16923 5412 16927 5468
rect 16927 5412 16983 5468
rect 16983 5412 16987 5468
rect 16923 5408 16987 5412
rect 2918 4924 2982 4928
rect 2918 4868 2922 4924
rect 2922 4868 2978 4924
rect 2978 4868 2982 4924
rect 2918 4864 2982 4868
rect 2998 4924 3062 4928
rect 2998 4868 3002 4924
rect 3002 4868 3058 4924
rect 3058 4868 3062 4924
rect 2998 4864 3062 4868
rect 3078 4924 3142 4928
rect 3078 4868 3082 4924
rect 3082 4868 3138 4924
rect 3138 4868 3142 4924
rect 3078 4864 3142 4868
rect 3158 4924 3222 4928
rect 3158 4868 3162 4924
rect 3162 4868 3218 4924
rect 3218 4868 3222 4924
rect 3158 4864 3222 4868
rect 6851 4924 6915 4928
rect 6851 4868 6855 4924
rect 6855 4868 6911 4924
rect 6911 4868 6915 4924
rect 6851 4864 6915 4868
rect 6931 4924 6995 4928
rect 6931 4868 6935 4924
rect 6935 4868 6991 4924
rect 6991 4868 6995 4924
rect 6931 4864 6995 4868
rect 7011 4924 7075 4928
rect 7011 4868 7015 4924
rect 7015 4868 7071 4924
rect 7071 4868 7075 4924
rect 7011 4864 7075 4868
rect 7091 4924 7155 4928
rect 7091 4868 7095 4924
rect 7095 4868 7151 4924
rect 7151 4868 7155 4924
rect 7091 4864 7155 4868
rect 10784 4924 10848 4928
rect 10784 4868 10788 4924
rect 10788 4868 10844 4924
rect 10844 4868 10848 4924
rect 10784 4864 10848 4868
rect 10864 4924 10928 4928
rect 10864 4868 10868 4924
rect 10868 4868 10924 4924
rect 10924 4868 10928 4924
rect 10864 4864 10928 4868
rect 10944 4924 11008 4928
rect 10944 4868 10948 4924
rect 10948 4868 11004 4924
rect 11004 4868 11008 4924
rect 10944 4864 11008 4868
rect 11024 4924 11088 4928
rect 11024 4868 11028 4924
rect 11028 4868 11084 4924
rect 11084 4868 11088 4924
rect 11024 4864 11088 4868
rect 14717 4924 14781 4928
rect 14717 4868 14721 4924
rect 14721 4868 14777 4924
rect 14777 4868 14781 4924
rect 14717 4864 14781 4868
rect 14797 4924 14861 4928
rect 14797 4868 14801 4924
rect 14801 4868 14857 4924
rect 14857 4868 14861 4924
rect 14797 4864 14861 4868
rect 14877 4924 14941 4928
rect 14877 4868 14881 4924
rect 14881 4868 14937 4924
rect 14937 4868 14941 4924
rect 14877 4864 14941 4868
rect 14957 4924 15021 4928
rect 14957 4868 14961 4924
rect 14961 4868 15017 4924
rect 15017 4868 15021 4924
rect 14957 4864 15021 4868
rect 4884 4380 4948 4384
rect 4884 4324 4888 4380
rect 4888 4324 4944 4380
rect 4944 4324 4948 4380
rect 4884 4320 4948 4324
rect 4964 4380 5028 4384
rect 4964 4324 4968 4380
rect 4968 4324 5024 4380
rect 5024 4324 5028 4380
rect 4964 4320 5028 4324
rect 5044 4380 5108 4384
rect 5044 4324 5048 4380
rect 5048 4324 5104 4380
rect 5104 4324 5108 4380
rect 5044 4320 5108 4324
rect 5124 4380 5188 4384
rect 5124 4324 5128 4380
rect 5128 4324 5184 4380
rect 5184 4324 5188 4380
rect 5124 4320 5188 4324
rect 8817 4380 8881 4384
rect 8817 4324 8821 4380
rect 8821 4324 8877 4380
rect 8877 4324 8881 4380
rect 8817 4320 8881 4324
rect 8897 4380 8961 4384
rect 8897 4324 8901 4380
rect 8901 4324 8957 4380
rect 8957 4324 8961 4380
rect 8897 4320 8961 4324
rect 8977 4380 9041 4384
rect 8977 4324 8981 4380
rect 8981 4324 9037 4380
rect 9037 4324 9041 4380
rect 8977 4320 9041 4324
rect 9057 4380 9121 4384
rect 9057 4324 9061 4380
rect 9061 4324 9117 4380
rect 9117 4324 9121 4380
rect 9057 4320 9121 4324
rect 12750 4380 12814 4384
rect 12750 4324 12754 4380
rect 12754 4324 12810 4380
rect 12810 4324 12814 4380
rect 12750 4320 12814 4324
rect 12830 4380 12894 4384
rect 12830 4324 12834 4380
rect 12834 4324 12890 4380
rect 12890 4324 12894 4380
rect 12830 4320 12894 4324
rect 12910 4380 12974 4384
rect 12910 4324 12914 4380
rect 12914 4324 12970 4380
rect 12970 4324 12974 4380
rect 12910 4320 12974 4324
rect 12990 4380 13054 4384
rect 12990 4324 12994 4380
rect 12994 4324 13050 4380
rect 13050 4324 13054 4380
rect 12990 4320 13054 4324
rect 16683 4380 16747 4384
rect 16683 4324 16687 4380
rect 16687 4324 16743 4380
rect 16743 4324 16747 4380
rect 16683 4320 16747 4324
rect 16763 4380 16827 4384
rect 16763 4324 16767 4380
rect 16767 4324 16823 4380
rect 16823 4324 16827 4380
rect 16763 4320 16827 4324
rect 16843 4380 16907 4384
rect 16843 4324 16847 4380
rect 16847 4324 16903 4380
rect 16903 4324 16907 4380
rect 16843 4320 16907 4324
rect 16923 4380 16987 4384
rect 16923 4324 16927 4380
rect 16927 4324 16983 4380
rect 16983 4324 16987 4380
rect 16923 4320 16987 4324
rect 2918 3836 2982 3840
rect 2918 3780 2922 3836
rect 2922 3780 2978 3836
rect 2978 3780 2982 3836
rect 2918 3776 2982 3780
rect 2998 3836 3062 3840
rect 2998 3780 3002 3836
rect 3002 3780 3058 3836
rect 3058 3780 3062 3836
rect 2998 3776 3062 3780
rect 3078 3836 3142 3840
rect 3078 3780 3082 3836
rect 3082 3780 3138 3836
rect 3138 3780 3142 3836
rect 3078 3776 3142 3780
rect 3158 3836 3222 3840
rect 3158 3780 3162 3836
rect 3162 3780 3218 3836
rect 3218 3780 3222 3836
rect 3158 3776 3222 3780
rect 6851 3836 6915 3840
rect 6851 3780 6855 3836
rect 6855 3780 6911 3836
rect 6911 3780 6915 3836
rect 6851 3776 6915 3780
rect 6931 3836 6995 3840
rect 6931 3780 6935 3836
rect 6935 3780 6991 3836
rect 6991 3780 6995 3836
rect 6931 3776 6995 3780
rect 7011 3836 7075 3840
rect 7011 3780 7015 3836
rect 7015 3780 7071 3836
rect 7071 3780 7075 3836
rect 7011 3776 7075 3780
rect 7091 3836 7155 3840
rect 7091 3780 7095 3836
rect 7095 3780 7151 3836
rect 7151 3780 7155 3836
rect 7091 3776 7155 3780
rect 10784 3836 10848 3840
rect 10784 3780 10788 3836
rect 10788 3780 10844 3836
rect 10844 3780 10848 3836
rect 10784 3776 10848 3780
rect 10864 3836 10928 3840
rect 10864 3780 10868 3836
rect 10868 3780 10924 3836
rect 10924 3780 10928 3836
rect 10864 3776 10928 3780
rect 10944 3836 11008 3840
rect 10944 3780 10948 3836
rect 10948 3780 11004 3836
rect 11004 3780 11008 3836
rect 10944 3776 11008 3780
rect 11024 3836 11088 3840
rect 11024 3780 11028 3836
rect 11028 3780 11084 3836
rect 11084 3780 11088 3836
rect 11024 3776 11088 3780
rect 14717 3836 14781 3840
rect 14717 3780 14721 3836
rect 14721 3780 14777 3836
rect 14777 3780 14781 3836
rect 14717 3776 14781 3780
rect 14797 3836 14861 3840
rect 14797 3780 14801 3836
rect 14801 3780 14857 3836
rect 14857 3780 14861 3836
rect 14797 3776 14861 3780
rect 14877 3836 14941 3840
rect 14877 3780 14881 3836
rect 14881 3780 14937 3836
rect 14937 3780 14941 3836
rect 14877 3776 14941 3780
rect 14957 3836 15021 3840
rect 14957 3780 14961 3836
rect 14961 3780 15017 3836
rect 15017 3780 15021 3836
rect 14957 3776 15021 3780
rect 4884 3292 4948 3296
rect 4884 3236 4888 3292
rect 4888 3236 4944 3292
rect 4944 3236 4948 3292
rect 4884 3232 4948 3236
rect 4964 3292 5028 3296
rect 4964 3236 4968 3292
rect 4968 3236 5024 3292
rect 5024 3236 5028 3292
rect 4964 3232 5028 3236
rect 5044 3292 5108 3296
rect 5044 3236 5048 3292
rect 5048 3236 5104 3292
rect 5104 3236 5108 3292
rect 5044 3232 5108 3236
rect 5124 3292 5188 3296
rect 5124 3236 5128 3292
rect 5128 3236 5184 3292
rect 5184 3236 5188 3292
rect 5124 3232 5188 3236
rect 8817 3292 8881 3296
rect 8817 3236 8821 3292
rect 8821 3236 8877 3292
rect 8877 3236 8881 3292
rect 8817 3232 8881 3236
rect 8897 3292 8961 3296
rect 8897 3236 8901 3292
rect 8901 3236 8957 3292
rect 8957 3236 8961 3292
rect 8897 3232 8961 3236
rect 8977 3292 9041 3296
rect 8977 3236 8981 3292
rect 8981 3236 9037 3292
rect 9037 3236 9041 3292
rect 8977 3232 9041 3236
rect 9057 3292 9121 3296
rect 9057 3236 9061 3292
rect 9061 3236 9117 3292
rect 9117 3236 9121 3292
rect 9057 3232 9121 3236
rect 12750 3292 12814 3296
rect 12750 3236 12754 3292
rect 12754 3236 12810 3292
rect 12810 3236 12814 3292
rect 12750 3232 12814 3236
rect 12830 3292 12894 3296
rect 12830 3236 12834 3292
rect 12834 3236 12890 3292
rect 12890 3236 12894 3292
rect 12830 3232 12894 3236
rect 12910 3292 12974 3296
rect 12910 3236 12914 3292
rect 12914 3236 12970 3292
rect 12970 3236 12974 3292
rect 12910 3232 12974 3236
rect 12990 3292 13054 3296
rect 12990 3236 12994 3292
rect 12994 3236 13050 3292
rect 13050 3236 13054 3292
rect 12990 3232 13054 3236
rect 16683 3292 16747 3296
rect 16683 3236 16687 3292
rect 16687 3236 16743 3292
rect 16743 3236 16747 3292
rect 16683 3232 16747 3236
rect 16763 3292 16827 3296
rect 16763 3236 16767 3292
rect 16767 3236 16823 3292
rect 16823 3236 16827 3292
rect 16763 3232 16827 3236
rect 16843 3292 16907 3296
rect 16843 3236 16847 3292
rect 16847 3236 16903 3292
rect 16903 3236 16907 3292
rect 16843 3232 16907 3236
rect 16923 3292 16987 3296
rect 16923 3236 16927 3292
rect 16927 3236 16983 3292
rect 16983 3236 16987 3292
rect 16923 3232 16987 3236
rect 2918 2748 2982 2752
rect 2918 2692 2922 2748
rect 2922 2692 2978 2748
rect 2978 2692 2982 2748
rect 2918 2688 2982 2692
rect 2998 2748 3062 2752
rect 2998 2692 3002 2748
rect 3002 2692 3058 2748
rect 3058 2692 3062 2748
rect 2998 2688 3062 2692
rect 3078 2748 3142 2752
rect 3078 2692 3082 2748
rect 3082 2692 3138 2748
rect 3138 2692 3142 2748
rect 3078 2688 3142 2692
rect 3158 2748 3222 2752
rect 3158 2692 3162 2748
rect 3162 2692 3218 2748
rect 3218 2692 3222 2748
rect 3158 2688 3222 2692
rect 6851 2748 6915 2752
rect 6851 2692 6855 2748
rect 6855 2692 6911 2748
rect 6911 2692 6915 2748
rect 6851 2688 6915 2692
rect 6931 2748 6995 2752
rect 6931 2692 6935 2748
rect 6935 2692 6991 2748
rect 6991 2692 6995 2748
rect 6931 2688 6995 2692
rect 7011 2748 7075 2752
rect 7011 2692 7015 2748
rect 7015 2692 7071 2748
rect 7071 2692 7075 2748
rect 7011 2688 7075 2692
rect 7091 2748 7155 2752
rect 7091 2692 7095 2748
rect 7095 2692 7151 2748
rect 7151 2692 7155 2748
rect 7091 2688 7155 2692
rect 10784 2748 10848 2752
rect 10784 2692 10788 2748
rect 10788 2692 10844 2748
rect 10844 2692 10848 2748
rect 10784 2688 10848 2692
rect 10864 2748 10928 2752
rect 10864 2692 10868 2748
rect 10868 2692 10924 2748
rect 10924 2692 10928 2748
rect 10864 2688 10928 2692
rect 10944 2748 11008 2752
rect 10944 2692 10948 2748
rect 10948 2692 11004 2748
rect 11004 2692 11008 2748
rect 10944 2688 11008 2692
rect 11024 2748 11088 2752
rect 11024 2692 11028 2748
rect 11028 2692 11084 2748
rect 11084 2692 11088 2748
rect 11024 2688 11088 2692
rect 14717 2748 14781 2752
rect 14717 2692 14721 2748
rect 14721 2692 14777 2748
rect 14777 2692 14781 2748
rect 14717 2688 14781 2692
rect 14797 2748 14861 2752
rect 14797 2692 14801 2748
rect 14801 2692 14857 2748
rect 14857 2692 14861 2748
rect 14797 2688 14861 2692
rect 14877 2748 14941 2752
rect 14877 2692 14881 2748
rect 14881 2692 14937 2748
rect 14937 2692 14941 2748
rect 14877 2688 14941 2692
rect 14957 2748 15021 2752
rect 14957 2692 14961 2748
rect 14961 2692 15017 2748
rect 15017 2692 15021 2748
rect 14957 2688 15021 2692
rect 4884 2204 4948 2208
rect 4884 2148 4888 2204
rect 4888 2148 4944 2204
rect 4944 2148 4948 2204
rect 4884 2144 4948 2148
rect 4964 2204 5028 2208
rect 4964 2148 4968 2204
rect 4968 2148 5024 2204
rect 5024 2148 5028 2204
rect 4964 2144 5028 2148
rect 5044 2204 5108 2208
rect 5044 2148 5048 2204
rect 5048 2148 5104 2204
rect 5104 2148 5108 2204
rect 5044 2144 5108 2148
rect 5124 2204 5188 2208
rect 5124 2148 5128 2204
rect 5128 2148 5184 2204
rect 5184 2148 5188 2204
rect 5124 2144 5188 2148
rect 8817 2204 8881 2208
rect 8817 2148 8821 2204
rect 8821 2148 8877 2204
rect 8877 2148 8881 2204
rect 8817 2144 8881 2148
rect 8897 2204 8961 2208
rect 8897 2148 8901 2204
rect 8901 2148 8957 2204
rect 8957 2148 8961 2204
rect 8897 2144 8961 2148
rect 8977 2204 9041 2208
rect 8977 2148 8981 2204
rect 8981 2148 9037 2204
rect 9037 2148 9041 2204
rect 8977 2144 9041 2148
rect 9057 2204 9121 2208
rect 9057 2148 9061 2204
rect 9061 2148 9117 2204
rect 9117 2148 9121 2204
rect 9057 2144 9121 2148
rect 12750 2204 12814 2208
rect 12750 2148 12754 2204
rect 12754 2148 12810 2204
rect 12810 2148 12814 2204
rect 12750 2144 12814 2148
rect 12830 2204 12894 2208
rect 12830 2148 12834 2204
rect 12834 2148 12890 2204
rect 12890 2148 12894 2204
rect 12830 2144 12894 2148
rect 12910 2204 12974 2208
rect 12910 2148 12914 2204
rect 12914 2148 12970 2204
rect 12970 2148 12974 2204
rect 12910 2144 12974 2148
rect 12990 2204 13054 2208
rect 12990 2148 12994 2204
rect 12994 2148 13050 2204
rect 13050 2148 13054 2204
rect 12990 2144 13054 2148
rect 16683 2204 16747 2208
rect 16683 2148 16687 2204
rect 16687 2148 16743 2204
rect 16743 2148 16747 2204
rect 16683 2144 16747 2148
rect 16763 2204 16827 2208
rect 16763 2148 16767 2204
rect 16767 2148 16823 2204
rect 16823 2148 16827 2204
rect 16763 2144 16827 2148
rect 16843 2204 16907 2208
rect 16843 2148 16847 2204
rect 16847 2148 16903 2204
rect 16903 2148 16907 2204
rect 16843 2144 16907 2148
rect 16923 2204 16987 2208
rect 16923 2148 16927 2204
rect 16927 2148 16983 2204
rect 16983 2148 16987 2204
rect 16923 2144 16987 2148
<< metal4 >>
rect 2910 15808 3230 15824
rect 2910 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3230 15808
rect 2910 14720 3230 15744
rect 2910 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3230 14720
rect 2910 13632 3230 14656
rect 2910 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3230 13632
rect 2910 12544 3230 13568
rect 2910 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3230 12544
rect 2910 11456 3230 12480
rect 2910 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3230 11456
rect 2910 10368 3230 11392
rect 2910 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3230 10368
rect 2910 9280 3230 10304
rect 2910 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3230 9280
rect 2910 8192 3230 9216
rect 2910 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3230 8192
rect 2910 7104 3230 8128
rect 2910 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3230 7104
rect 2910 6016 3230 7040
rect 2910 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3230 6016
rect 2910 4928 3230 5952
rect 2910 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3230 4928
rect 2910 3840 3230 4864
rect 2910 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3230 3840
rect 2910 2752 3230 3776
rect 2910 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3230 2752
rect 2910 2128 3230 2688
rect 4876 15264 5196 15824
rect 4876 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5196 15264
rect 4876 14176 5196 15200
rect 4876 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5196 14176
rect 4876 13088 5196 14112
rect 4876 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5196 13088
rect 4876 12000 5196 13024
rect 4876 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5196 12000
rect 4876 10912 5196 11936
rect 4876 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5196 10912
rect 4876 9824 5196 10848
rect 4876 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5196 9824
rect 4876 8736 5196 9760
rect 4876 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5196 8736
rect 4876 7648 5196 8672
rect 4876 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5196 7648
rect 4876 6560 5196 7584
rect 4876 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5196 6560
rect 4876 5472 5196 6496
rect 4876 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5196 5472
rect 4876 4384 5196 5408
rect 4876 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5196 4384
rect 4876 3296 5196 4320
rect 4876 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5196 3296
rect 4876 2208 5196 3232
rect 4876 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5196 2208
rect 4876 2128 5196 2144
rect 6843 15808 7163 15824
rect 6843 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7163 15808
rect 6843 14720 7163 15744
rect 6843 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7163 14720
rect 6843 13632 7163 14656
rect 6843 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7163 13632
rect 6843 12544 7163 13568
rect 6843 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7163 12544
rect 6843 11456 7163 12480
rect 6843 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7163 11456
rect 6843 10368 7163 11392
rect 6843 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7163 10368
rect 6843 9280 7163 10304
rect 6843 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7163 9280
rect 6843 8192 7163 9216
rect 6843 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7163 8192
rect 6843 7104 7163 8128
rect 6843 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7163 7104
rect 6843 6016 7163 7040
rect 6843 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7163 6016
rect 6843 4928 7163 5952
rect 6843 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7163 4928
rect 6843 3840 7163 4864
rect 6843 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7163 3840
rect 6843 2752 7163 3776
rect 6843 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7163 2752
rect 6843 2128 7163 2688
rect 8809 15264 9129 15824
rect 8809 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9129 15264
rect 8809 14176 9129 15200
rect 8809 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9129 14176
rect 8809 13088 9129 14112
rect 8809 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9129 13088
rect 8809 12000 9129 13024
rect 8809 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9129 12000
rect 8809 10912 9129 11936
rect 8809 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9129 10912
rect 8809 9824 9129 10848
rect 8809 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9129 9824
rect 8809 8736 9129 9760
rect 8809 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9129 8736
rect 8809 7648 9129 8672
rect 8809 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9129 7648
rect 8809 6560 9129 7584
rect 8809 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9129 6560
rect 8809 5472 9129 6496
rect 8809 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9129 5472
rect 8809 4384 9129 5408
rect 8809 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9129 4384
rect 8809 3296 9129 4320
rect 8809 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9129 3296
rect 8809 2208 9129 3232
rect 8809 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9129 2208
rect 8809 2128 9129 2144
rect 10776 15808 11096 15824
rect 10776 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11096 15808
rect 10776 14720 11096 15744
rect 10776 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11096 14720
rect 10776 13632 11096 14656
rect 10776 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11096 13632
rect 10776 12544 11096 13568
rect 10776 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11096 12544
rect 10776 11456 11096 12480
rect 10776 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11096 11456
rect 10776 10368 11096 11392
rect 10776 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11096 10368
rect 10776 9280 11096 10304
rect 10776 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11096 9280
rect 10776 8192 11096 9216
rect 10776 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11096 8192
rect 10776 7104 11096 8128
rect 10776 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11096 7104
rect 10776 6016 11096 7040
rect 10776 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11096 6016
rect 10776 4928 11096 5952
rect 10776 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11096 4928
rect 10776 3840 11096 4864
rect 10776 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11096 3840
rect 10776 2752 11096 3776
rect 10776 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11096 2752
rect 10776 2128 11096 2688
rect 12742 15264 13062 15824
rect 12742 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13062 15264
rect 12742 14176 13062 15200
rect 12742 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13062 14176
rect 12742 13088 13062 14112
rect 12742 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13062 13088
rect 12742 12000 13062 13024
rect 12742 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13062 12000
rect 12742 10912 13062 11936
rect 12742 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13062 10912
rect 12742 9824 13062 10848
rect 12742 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13062 9824
rect 12742 8736 13062 9760
rect 12742 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13062 8736
rect 12742 7648 13062 8672
rect 12742 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13062 7648
rect 12742 6560 13062 7584
rect 12742 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13062 6560
rect 12742 5472 13062 6496
rect 12742 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13062 5472
rect 12742 4384 13062 5408
rect 12742 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13062 4384
rect 12742 3296 13062 4320
rect 12742 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13062 3296
rect 12742 2208 13062 3232
rect 12742 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13062 2208
rect 12742 2128 13062 2144
rect 14709 15808 15029 15824
rect 14709 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15029 15808
rect 14709 14720 15029 15744
rect 14709 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15029 14720
rect 14709 13632 15029 14656
rect 14709 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15029 13632
rect 14709 12544 15029 13568
rect 14709 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15029 12544
rect 14709 11456 15029 12480
rect 14709 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15029 11456
rect 14709 10368 15029 11392
rect 14709 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15029 10368
rect 14709 9280 15029 10304
rect 14709 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15029 9280
rect 14709 8192 15029 9216
rect 14709 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15029 8192
rect 14709 7104 15029 8128
rect 14709 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15029 7104
rect 14709 6016 15029 7040
rect 14709 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15029 6016
rect 14709 4928 15029 5952
rect 14709 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15029 4928
rect 14709 3840 15029 4864
rect 14709 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15029 3840
rect 14709 2752 15029 3776
rect 14709 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15029 2752
rect 14709 2128 15029 2688
rect 16675 15264 16995 15824
rect 16675 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16995 15264
rect 16675 14176 16995 15200
rect 16675 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16995 14176
rect 16675 13088 16995 14112
rect 16675 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16995 13088
rect 16675 12000 16995 13024
rect 16675 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16995 12000
rect 16675 10912 16995 11936
rect 16675 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16995 10912
rect 16675 9824 16995 10848
rect 16675 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16995 9824
rect 16675 8736 16995 9760
rect 16675 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16995 8736
rect 16675 7648 16995 8672
rect 16675 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16995 7648
rect 16675 6560 16995 7584
rect 16675 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16995 6560
rect 16675 5472 16995 6496
rect 16675 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16995 5472
rect 16675 4384 16995 5408
rect 16675 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16995 4384
rect 16675 3296 16995 4320
rect 16675 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16995 3296
rect 16675 2208 16995 3232
rect 16675 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16995 2208
rect 16675 2128 16995 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__59__C dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 10580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_reg_clk_A
timestamp 1673029049
transform -1 0 14444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1673029049
transform -1 0 5428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1673029049
transform -1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1673029049
transform -1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1673029049
transform -1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1673029049
transform -1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1673029049
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1673029049
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47
timestamp 1673029049
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1673029049
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1673029049
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1673029049
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1673029049
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1673029049
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1673029049
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1673029049
transform 1 0 9752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1673029049
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1673029049
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1673029049
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1673029049
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1673029049
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1673029049
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1673029049
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1673029049
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1673029049
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1673029049
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1673029049
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1673029049
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1673029049
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1673029049
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1673029049
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp 1673029049
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_80
timestamp 1673029049
transform 1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_88
timestamp 1673029049
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1673029049
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1673029049
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1673029049
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1673029049
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_138
timestamp 1673029049
transform 1 0 13800 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1673029049
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1673029049
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1673029049
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1673029049
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1673029049
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1673029049
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1673029049
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1673029049
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1673029049
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1673029049
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1673029049
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1673029049
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1673029049
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1673029049
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1673029049
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_125
timestamp 1673029049
transform 1 0 12604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1673029049
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1673029049
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 1673029049
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1673029049
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1673029049
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1673029049
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1673029049
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1673029049
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1673029049
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1673029049
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1673029049
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1673029049
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1673029049
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_82
timestamp 1673029049
transform 1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_91
timestamp 1673029049
transform 1 0 9476 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1673029049
transform 1 0 10212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1673029049
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1673029049
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1673029049
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1673029049
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1673029049
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_134
timestamp 1673029049
transform 1 0 13432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_140
timestamp 1673029049
transform 1 0 13984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_146
timestamp 1673029049
transform 1 0 14536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1673029049
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1673029049
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1673029049
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1673029049
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1673029049
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1673029049
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1673029049
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1673029049
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1673029049
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1673029049
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1673029049
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_107
timestamp 1673029049
transform 1 0 10948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1673029049
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_125
timestamp 1673029049
transform 1 0 12604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1673029049
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1673029049
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_155
timestamp 1673029049
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_162
timestamp 1673029049
transform 1 0 16008 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1673029049
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1673029049
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1673029049
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1673029049
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1673029049
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1673029049
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1673029049
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp 1673029049
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_77
timestamp 1673029049
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_92
timestamp 1673029049
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1673029049
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1673029049
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_120
timestamp 1673029049
transform 1 0 12144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_129
timestamp 1673029049
transform 1 0 12972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_138
timestamp 1673029049
transform 1 0 13800 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1673029049
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1673029049
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1673029049
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1673029049
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1673029049
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1673029049
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1673029049
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1673029049
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1673029049
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1673029049
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1673029049
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1673029049
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp 1673029049
transform 1 0 10764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_112
timestamp 1673029049
transform 1 0 11408 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1673029049
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1673029049
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1673029049
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1673029049
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1673029049
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1673029049
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1673029049
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1673029049
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1673029049
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1673029049
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1673029049
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1673029049
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1673029049
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1673029049
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_81
timestamp 1673029049
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1673029049
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_94
timestamp 1673029049
transform 1 0 9752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1673029049
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1673029049
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1673029049
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1673029049
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_131
timestamp 1673029049
transform 1 0 13156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_144
timestamp 1673029049
transform 1 0 14352 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_156
timestamp 1673029049
transform 1 0 15456 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1673029049
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1673029049
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1673029049
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1673029049
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1673029049
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1673029049
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1673029049
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1673029049
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1673029049
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1673029049
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1673029049
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_101
timestamp 1673029049
transform 1 0 10396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_113
timestamp 1673029049
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1673029049
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1673029049
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1673029049
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp 1673029049
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1673029049
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1673029049
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1673029049
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1673029049
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1673029049
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1673029049
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1673029049
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1673029049
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1673029049
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1673029049
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1673029049
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1673029049
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1673029049
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1673029049
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1673029049
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1673029049
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1673029049
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1673029049
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1673029049
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1673029049
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1673029049
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1673029049
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1673029049
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1673029049
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1673029049
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1673029049
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1673029049
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1673029049
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1673029049
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1673029049
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1673029049
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1673029049
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1673029049
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1673029049
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1673029049
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp 1673029049
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1673029049
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1673029049
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1673029049
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1673029049
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1673029049
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1673029049
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1673029049
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1673029049
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1673029049
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1673029049
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1673029049
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1673029049
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1673029049
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1673029049
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1673029049
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1673029049
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1673029049
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1673029049
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1673029049
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1673029049
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1673029049
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1673029049
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1673029049
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1673029049
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1673029049
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1673029049
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1673029049
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1673029049
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1673029049
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1673029049
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1673029049
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1673029049
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1673029049
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1673029049
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1673029049
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_165
timestamp 1673029049
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1673029049
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1673029049
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1673029049
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1673029049
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1673029049
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1673029049
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1673029049
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1673029049
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1673029049
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1673029049
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1673029049
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1673029049
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1673029049
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1673029049
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1673029049
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1673029049
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1673029049
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1673029049
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1673029049
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1673029049
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1673029049
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1673029049
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1673029049
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1673029049
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1673029049
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1673029049
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1673029049
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1673029049
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1673029049
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1673029049
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1673029049
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1673029049
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1673029049
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1673029049
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1673029049
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_165
timestamp 1673029049
transform 1 0 16284 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1673029049
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1673029049
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1673029049
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1673029049
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1673029049
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1673029049
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1673029049
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1673029049
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1673029049
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1673029049
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1673029049
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1673029049
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1673029049
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1673029049
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1673029049
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1673029049
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1673029049
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1673029049
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1673029049
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1673029049
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1673029049
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1673029049
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1673029049
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1673029049
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1673029049
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1673029049
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1673029049
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1673029049
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1673029049
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1673029049
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1673029049
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1673029049
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1673029049
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1673029049
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1673029049
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_165
timestamp 1673029049
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1673029049
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1673029049
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1673029049
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1673029049
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1673029049
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1673029049
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1673029049
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1673029049
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1673029049
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1673029049
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1673029049
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1673029049
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1673029049
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1673029049
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1673029049
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1673029049
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1673029049
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1673029049
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1673029049
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1673029049
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1673029049
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1673029049
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1673029049
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1673029049
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1673029049
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1673029049
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1673029049
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1673029049
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1673029049
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1673029049
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1673029049
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1673029049
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1673029049
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1673029049
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1673029049
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_165
timestamp 1673029049
transform 1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1673029049
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1673029049
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1673029049
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1673029049
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1673029049
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1673029049
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1673029049
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1673029049
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1673029049
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1673029049
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1673029049
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1673029049
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1673029049
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1673029049
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1673029049
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1673029049
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1673029049
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1673029049
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1673029049
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1673029049
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1673029049
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1673029049
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1673029049
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1673029049
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1673029049
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1673029049
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1673029049
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1673029049
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1673029049
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1673029049
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1673029049
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1673029049
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1673029049
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1673029049
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1673029049
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1673029049
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1673029049
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1673029049
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1673029049
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1673029049
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1673029049
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1673029049
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1673029049
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1673029049
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1673029049
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1673029049
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1673029049
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1673029049
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1673029049
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1673029049
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1673029049
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1673029049
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1673029049
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1673029049
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1673029049
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1673029049
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1673029049
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1673029049
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1673029049
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1673029049
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1673029049
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1673029049
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1673029049
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1673029049
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1673029049
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1673029049
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1673029049
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1673029049
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1673029049
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1673029049
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1673029049
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1673029049
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1673029049
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1673029049
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1673029049
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1673029049
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1673029049
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1673029049
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1673029049
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1673029049
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1673029049
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1673029049
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1673029049
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1673029049
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1673029049
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1673029049
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1673029049
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1673029049
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1673029049
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1673029049
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1673029049
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_9
timestamp 1673029049
transform 1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1673029049
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1673029049
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1673029049
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_35
timestamp 1673029049
transform 1 0 4324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_47
timestamp 1673029049
transform 1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_54
timestamp 1673029049
transform 1 0 6072 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_57
timestamp 1673029049
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1673029049
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_73
timestamp 1673029049
transform 1 0 7820 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_78
timestamp 1673029049
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1673029049
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1673029049
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1673029049
transform 1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1673029049
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_113
timestamp 1673029049
transform 1 0 11500 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1673029049
transform 1 0 12236 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_126
timestamp 1673029049
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1673029049
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1673029049
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1673029049
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_150
timestamp 1673029049
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_166
timestamp 1673029049
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1673029049
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1673029049
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1673029049
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1673029049
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1673029049
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1673029049
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1673029049
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1673029049
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1673029049
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1673029049
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1673029049
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1673029049
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1673029049
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1673029049
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1673029049
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1673029049
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1673029049
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1673029049
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1673029049
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1673029049
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1673029049
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1673029049
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1673029049
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1673029049
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1673029049
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1673029049
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1673029049
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1673029049
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1673029049
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1673029049
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1673029049
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1673029049
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1673029049
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1673029049
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1673029049
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1673029049
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1673029049
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1673029049
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1673029049
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1673029049
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1673029049
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1673029049
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1673029049
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1673029049
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1673029049
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1673029049
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1673029049
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1673029049
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1673029049
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1673029049
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1673029049
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1673029049
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1673029049
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1673029049
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1673029049
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1673029049
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1673029049
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1673029049
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1673029049
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1673029049
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1673029049
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1673029049
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1673029049
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1673029049
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1673029049
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1673029049
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1673029049
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1673029049
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1673029049
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1673029049
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1673029049
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1673029049
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1673029049
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1673029049
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1673029049
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1673029049
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1673029049
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1673029049
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1673029049
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1673029049
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1673029049
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1673029049
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1673029049
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1673029049
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1673029049
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1673029049
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1673029049
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1673029049
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1673029049
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1673029049
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1673029049
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1673029049
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or4b_2  _33_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _34_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12880 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _35_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 11776 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _36_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 10120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _37_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _38_
timestamp 1673029049
transform -1 0 9476 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1673029049
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _40_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 11040 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _41_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12144 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _42_
timestamp 1673029049
transform 1 0 12512 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1673029049
transform 1 0 12604 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _44_
timestamp 1673029049
transform 1 0 11960 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _45_
timestamp 1673029049
transform -1 0 12144 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1673029049
transform -1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _47_
timestamp 1673029049
transform 1 0 13340 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1673029049
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _49_
timestamp 1673029049
transform -1 0 13432 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1673029049
transform -1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _51_
timestamp 1673029049
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _52_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1673029049
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _54_
timestamp 1673029049
transform 1 0 11408 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1673029049
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _56_
timestamp 1673029049
transform -1 0 8648 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1673029049
transform -1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _58_
timestamp 1673029049
transform 1 0 9292 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _59_
timestamp 1673029049
transform -1 0 12236 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _60_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 10948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _61_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 14260 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _62_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 14536 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _63_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 10304 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _64_
timestamp 1673029049
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _65_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 13156 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlxtn_1  _66_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 9844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _67_
timestamp 1673029049
transform 1 0 9108 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _68_
timestamp 1673029049
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _69_
timestamp 1673029049
transform 1 0 11684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _70_
timestamp 1673029049
transform 1 0 13248 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _71_
timestamp 1673029049
transform 1 0 14260 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_4  _72_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 9384 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxtn_1  _73_
timestamp 1673029049
transform 1 0 11684 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _74_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 16376 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _75_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 13800 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _76_
timestamp 1673029049
transform -1 0 16376 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _77_
timestamp 1673029049
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_reg_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 16376 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_reg_clk
timestamp 1673029049
transform 1 0 14536 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_reg_clk
timestamp 1673029049
transform 1 0 14536 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1673029049
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1673029049
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1673029049
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1673029049
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1673029049
transform -1 0 4324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1673029049
transform -1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1673029049
transform -1 0 8280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1673029049
transform -1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1673029049
transform -1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1673029049
transform -1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1673029049
transform 1 0 16008 0 1 15232
box -38 -48 406 592
<< labels >>
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 reg_addr[0]
port 0 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 reg_addr[1]
port 1 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 reg_addr[2]
port 2 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 reg_bus
port 3 nsew signal bidirectional
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 reg_clk
port 4 nsew signal input
flabel metal2 s 1214 17200 1270 18000 0 FreeSans 224 90 0 0 reg_data[0]
port 5 nsew signal tristate
flabel metal2 s 3422 17200 3478 18000 0 FreeSans 224 90 0 0 reg_data[1]
port 6 nsew signal tristate
flabel metal2 s 5630 17200 5686 18000 0 FreeSans 224 90 0 0 reg_data[2]
port 7 nsew signal tristate
flabel metal2 s 7838 17200 7894 18000 0 FreeSans 224 90 0 0 reg_data[3]
port 8 nsew signal tristate
flabel metal2 s 10046 17200 10102 18000 0 FreeSans 224 90 0 0 reg_data[4]
port 9 nsew signal tristate
flabel metal2 s 12254 17200 12310 18000 0 FreeSans 224 90 0 0 reg_data[5]
port 10 nsew signal tristate
flabel metal2 s 14462 17200 14518 18000 0 FreeSans 224 90 0 0 reg_data[6]
port 11 nsew signal tristate
flabel metal2 s 16670 17200 16726 18000 0 FreeSans 224 90 0 0 reg_data[7]
port 12 nsew signal tristate
flabel metal2 s 1582 0 1638 800 0 FreeSans 224 90 0 0 reg_dir
port 13 nsew signal input
flabel metal4 s 2910 2128 3230 15824 0 FreeSans 1920 90 0 0 vcc
port 14 nsew power bidirectional
flabel metal4 s 6843 2128 7163 15824 0 FreeSans 1920 90 0 0 vcc
port 14 nsew power bidirectional
flabel metal4 s 10776 2128 11096 15824 0 FreeSans 1920 90 0 0 vcc
port 14 nsew power bidirectional
flabel metal4 s 14709 2128 15029 15824 0 FreeSans 1920 90 0 0 vcc
port 14 nsew power bidirectional
flabel metal4 s 4876 2128 5196 15824 0 FreeSans 1920 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 8809 2128 9129 15824 0 FreeSans 1920 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 12742 2128 13062 15824 0 FreeSans 1920 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 16675 2128 16995 15824 0 FreeSans 1920 90 0 0 vss
port 15 nsew ground bidirectional
rlabel metal1 8970 15776 8970 15776 0 vcc
rlabel via1 9049 15232 9049 15232 0 vss
rlabel metal1 9384 2618 9384 2618 0 _00_
rlabel metal2 11730 2788 11730 2788 0 _01_
rlabel metal1 8556 4250 8556 4250 0 _02_
rlabel metal1 10028 6630 10028 6630 0 _03_
rlabel metal2 9154 5916 9154 5916 0 _04_
rlabel metal2 12650 6324 12650 6324 0 _05_
rlabel metal2 11362 6052 11362 6052 0 _06_
rlabel metal2 13294 6052 13294 6052 0 _07_
rlabel metal1 13432 3706 13432 3706 0 _08_
rlabel via1 16058 3502 16058 3502 0 _09_
rlabel metal1 13344 2414 13344 2414 0 _10_
rlabel metal1 14628 3162 14628 3162 0 _11_
rlabel metal2 9246 3536 9246 3536 0 _12_
rlabel metal1 11730 4556 11730 4556 0 _13_
rlabel metal2 11362 5219 11362 5219 0 _14_
rlabel metal1 13248 4522 13248 4522 0 _15_
rlabel metal1 9062 4012 9062 4012 0 _16_
rlabel metal1 11270 4114 11270 4114 0 _17_
rlabel metal1 12558 5236 12558 5236 0 _18_
rlabel metal1 13018 5338 13018 5338 0 _19_
rlabel metal1 12604 3910 12604 3910 0 _20_
rlabel metal1 11454 5338 11454 5338 0 _21_
rlabel metal1 13616 5338 13616 5338 0 _22_
rlabel metal1 12512 3502 12512 3502 0 _23_
rlabel metal1 8786 2414 8786 2414 0 _24_
rlabel metal2 11914 2890 11914 2890 0 _25_
rlabel metal2 8418 4284 8418 4284 0 _26_
rlabel metal1 10166 4046 10166 4046 0 _27_
rlabel metal1 11086 4590 11086 4590 0 _28_
rlabel metal1 10350 4114 10350 4114 0 _29_
rlabel metal1 14812 4114 14812 4114 0 _30_
rlabel metal1 12466 4046 12466 4046 0 _31_
rlabel metal2 9706 3468 9706 3468 0 _32_
rlabel metal2 14582 4148 14582 4148 0 clknet_0_reg_clk
rlabel metal1 15870 2516 15870 2516 0 clknet_1_0__leaf_reg_clk
rlabel metal2 16330 4624 16330 4624 0 clknet_1_1__leaf_reg_clk
rlabel metal1 4830 2312 4830 2312 0 net1
rlabel metal1 13156 6086 13156 6086 0 net10
rlabel metal1 14812 6086 14812 6086 0 net11
rlabel metal1 15272 4794 15272 4794 0 net12
rlabel metal1 8142 2346 8142 2346 0 net2
rlabel metal1 8280 2414 8280 2414 0 net3
rlabel metal2 8418 2822 8418 2822 0 net4
rlabel metal1 2116 15470 2116 15470 0 net5
rlabel metal2 4278 10404 4278 10404 0 net6
rlabel metal1 10672 6086 10672 6086 0 net7
rlabel metal1 10396 4658 10396 4658 0 net8
rlabel metal2 13662 6188 13662 6188 0 net9
rlabel metal1 4600 2414 4600 2414 0 reg_addr[0]
rlabel metal1 7406 2414 7406 2414 0 reg_addr[1]
rlabel metal1 10580 2414 10580 2414 0 reg_addr[2]
rlabel metal1 12190 3026 12190 3026 0 reg_bus
rlabel metal2 16330 1894 16330 1894 0 reg_clk
rlabel metal1 1472 15674 1472 15674 0 reg_data[0]
rlabel metal1 3772 15674 3772 15674 0 reg_data[1]
rlabel metal2 5757 17340 5757 17340 0 reg_data[2]
rlabel metal2 7965 17340 7965 17340 0 reg_data[3]
rlabel metal2 10173 17340 10173 17340 0 reg_data[4]
rlabel metal2 12335 17340 12335 17340 0 reg_data[5]
rlabel metal1 14582 15674 14582 15674 0 reg_data[6]
rlabel metal2 16698 16500 16698 16500 0 reg_data[7]
rlabel metal1 1656 2414 1656 2414 0 reg_dir
rlabel metal1 11500 3570 11500 3570 0 t\[0\]
rlabel metal1 13202 5134 13202 5134 0 t\[1\]
rlabel metal1 9016 4114 9016 4114 0 t\[2\]
<< properties >>
string FIXED_BBOX 0 0 18000 18000
<< end >>
