* NGSPICE file created from spi_device.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

.subckt spi_device reg_addr[0] reg_addr[1] reg_addr[2] reg_bus reg_clk reg_dir spi_clk
+ spi_miso spi_mosi spi_sel vcc vss
XFILLER_22_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_9_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_12_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_66_ _01_ _10_ vss vss vcc vcc net4 sky130_fd_sc_hd__dlxtn_1
XFILLER_2_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_2_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_49_ _26_ vss vss vcc vcc next_state\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_18_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_53 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_19_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_3 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_15_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
Xoutput7 net7 vss vss vcc vcc reg_dir sky130_fd_sc_hd__buf_2
XFILLER_16_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_112 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_9_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_12_11 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_65_ net2 vss vss vcc vcc _16_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f_spi_clk clknet_0_spi_clk vss vss vcc vcc clknet_1_1__leaf_spi_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_23_54 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_23_65 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_2_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_0_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_48_ pres_state\[1\] vss vss vcc vcc _26_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_16_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_16_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
Xoutput8 net8 vss vss vcc vcc spi_miso sky130_fd_sc_hd__buf_2
XFILLER_15_77 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_113 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_23 vss vss vcc vcc sky130_fd_sc_hd__decap_4
X_64_ net2 vss vss vcc vcc _15_ sky130_fd_sc_hd__inv_2
XFILLER_23_44 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_47_ _25_ vss vss vcc vcc next_state\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_9_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_15_34 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_89 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_114 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_63_ net2 vss vss vcc vcc _14_ sky130_fd_sc_hd__inv_2
XFILLER_23_78 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_9_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_46_ _17_ _24_ vss vss vcc vcc _25_ sky130_fd_sc_hd__or2b_1
XFILLER_18_34 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_1_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_57 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XTAP_115 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_62_ net2 vss vss vcc vcc _13_ sky130_fd_sc_hd__inv_2
XFILLER_23_57 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_9_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_45_ pres_state\[1\] net2 vss vss vcc vcc _24_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f_spi_clk clknet_0_spi_clk vss vss vcc vcc clknet_1_0__leaf_spi_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_1_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_58 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_20_25 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_19_110 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_6_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_15_14 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XTAP_116 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_61_ net2 vss vss vcc vcc _12_ sky130_fd_sc_hd__inv_2
XFILLER_0_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_44_ _17_ _23_ pres_state\[1\] vss vss vcc vcc _09_ sky130_fd_sc_hd__a21o_1
XFILLER_18_25 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_1_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_90 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_80 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XTAP_106 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_8_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_10_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_60_ _31_ vss vss vcc vcc _07_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_9_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_43_ t\[1\] t\[2\] t\[0\] vss vss vcc vcc _23_ sky130_fd_sc_hd__or3b_1
XFILLER_1_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_19_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_6_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_49 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XTAP_107 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_92 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_1 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_8_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_5_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_42_ _22_ vss vss vcc vcc _08_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_102 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_10_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XTAP_108 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_12_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_17 vss vss vcc vcc sky130_fd_sc_hd__decap_4
X_41_ pres_state\[1\] _21_ vss vss vcc vcc _22_ sky130_fd_sc_hd__or2_1
XFILLER_24_82 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_20_29 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_19_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_161 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XTAP_109 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_61 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_16_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_22_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_3 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_15_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_12_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_5_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_40_ t\[1\] t\[2\] t\[0\] pres_state\[0\] vss vss vcc vcc _21_ sky130_fd_sc_hd__o31a_1
XFILLER_18_29 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_spi_clk_A spi_clk vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_19_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_4 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_12_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_2_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_62 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_1_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_19_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_24_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_5 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_16_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_4_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_53 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_24_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_74 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_10_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_153 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_16_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_6 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_21_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_16_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_1_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_24_97 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_1_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
Xinput1 spi_mosi vss vss vcc vcc net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XTAP_90 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_54 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_21_43 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_21_21 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_7 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_23_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_21_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_54 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_7_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_4_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_1_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_13_11 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_13_33 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_54 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_24_10 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XANTENNA_input2_A spi_sel vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_1_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
Xinput2 spi_sel vss vss vcc vcc net2 sky130_fd_sc_hd__clkbuf_2
XTAP_80 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_166 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XPHY_8 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_21_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_66 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_44 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_4_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_1_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_23 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_13_45 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_24_33 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_1_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_92 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_66 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_18_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_101 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_9 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_101 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_15_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_21_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_104 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_16_78 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_4_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_1_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_1_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_77_ _01_ _09_ vss vss vcc vcc net3 sky130_fd_sc_hd__dlxtn_1
XTAP_93 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_78 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_12 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_18_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_18_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_68 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_57 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_21_13 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_7_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_4_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_13_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_1_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_57 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_24_24 vss vss vcc vcc sky130_fd_sc_hd__decap_4
X_76_ _01_ _08_ vss vss vcc vcc net7 sky130_fd_sc_hd__dlxtn_1
XFILLER_1_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_57 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XTAP_94 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_83 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_24_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_59_ _17_ vss vss vcc vcc _31_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_47 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_7_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_11_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_14_3 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_13_15 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_1_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_1_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_8_8 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_5_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_75_ _00_ _07_ vss vss vcc vcc net6 sky130_fd_sc_hd__dlxtn_1
XFILLER_19_36 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XTAP_95 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XTAP_84 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_137 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_2_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_58_ _30_ vss vss vcc vcc _01_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_26 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_16_15 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_7_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_4_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_96 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_74_ net1 _06_ vss vss vcc vcc reg_bus sky130_fd_sc_hd__dlxtn_2
XTAP_52 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_57_ pres_state\[1\] net1 pres_state\[0\] vss vss vcc vcc _30_ sky130_fd_sc_hd__and3b_1
XFILLER_11_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_24_38 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_5_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XTAP_97 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_73_ reg_bus _05_ vss vss vcc vcc net8 sky130_fd_sc_hd__dlxtn_1
XTAP_53 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_49 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_10_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_106 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_56_ _29_ vss vss vcc vcc _00_ sky130_fd_sc_hd__buf_1
XFILLER_2_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_16_9 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_39_ _17_ pres_state\[1\] net7 vss vss vcc vcc _06_ sky130_fd_sc_hd__nand3b_1
XFILLER_20_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_3 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_0_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_17 vss vss vcc vcc sky130_fd_sc_hd__decap_4
X_72_ clknet_1_0__leaf_spi_clk next_state\[1\] _16_ vss vss vcc vcc pres_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_98 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_50 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_72 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_55_ _17_ pres_state\[1\] clknet_1_0__leaf_spi_clk vss vss vcc vcc _29_ sky130_fd_sc_hd__and3b_2
XFILLER_2_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_20_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_20_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_29 vss vss vcc vcc sky130_fd_sc_hd__fill_2
X_38_ _20_ vss vss vcc vcc _05_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_3_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_0_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_29 vss vss vcc vcc sky130_fd_sc_hd__decap_4
X_71_ clknet_1_0__leaf_spi_clk next_state\[0\] _15_ vss vss vcc vcc pres_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_62 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XTAP_99 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_54_ _19_ _28_ _24_ _17_ vss vss vcc vcc _04_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_37_ pres_state\[0\] net7 pres_state\[1\] vss vss vcc vcc _20_ sky130_fd_sc_hd__or3b_1
XFILLER_16_19 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_7_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_0_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_14_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_70_ clknet_1_1__leaf_spi_clk _04_ _14_ vss vss vcc vcc t\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_56 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_40 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_53_ t\[1\] t\[0\] t\[2\] vss vss vcc vcc _28_ sky130_fd_sc_hd__a21bo_1
XFILLER_17_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_2_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_15_109 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_14_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_36_ _17_ _19_ pres_state\[1\] vss vss vcc vcc _11_ sky130_fd_sc_hd__a21o_1
XFILLER_22_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_52 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_7_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_7_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_9 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_63 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_41 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_5_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_10_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_57 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_52_ _17_ _24_ _27_ vss vss vcc vcc _03_ sky130_fd_sc_hd__o21a_1
XPHY_30 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_23_110 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_14_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_35_ t\[2\] t\[0\] t\[1\] vss vss vcc vcc _19_ sky130_fd_sc_hd__nand3b_1
XFILLER_14_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_11_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_4_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_75 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_12_7 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_14_21 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XTAP_58 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_20 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_31 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_51_ t\[1\] t\[0\] vss vss vcc vcc _27_ sky130_fd_sc_hd__xor2_1
XFILLER_11_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_34_ _17_ _18_ pres_state\[1\] vss vss vcc vcc _10_ sky130_fd_sc_hd__a21o_1
Xclkbuf_0_spi_clk spi_clk vss vss vcc vcc clknet_0_spi_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_14_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_0_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_11_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_59 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_18_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_32 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_10 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_21 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_50_ _17_ _24_ t\[0\] vss vss vcc vcc _02_ sky130_fd_sc_hd__o21ba_1
XFILLER_23_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_33_ t\[2\] t\[0\] t\[1\] vss vss vcc vcc _18_ sky130_fd_sc_hd__or3b_1
XFILLER_11_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_17_33 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_3_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_0_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_44 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_33 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_11 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_22 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_2_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_102 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_11_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_32_ pres_state\[0\] vss vss vcc vcc _17_ sky130_fd_sc_hd__buf_2
XFILLER_9_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_22_78 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_11_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_11_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_3 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_6_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_14 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_0_81 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_0_137 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_5_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_12 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_45 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_34 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_2_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_23 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_23_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_22_68 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_8_26 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_17_57 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_3_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_46 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_35 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_13 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_9_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_24 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_23_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_3_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_3 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_23_90 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_47 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_36 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_14 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_25 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_26 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_10_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_9_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_14_38 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_70 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_48 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_37 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_6_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_15 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_26 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_20_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_13_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_0_9 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_0_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_81 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_20_82 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XPHY_49 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_38 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_16 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_27 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_10_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_12_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_17_17 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_0_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_53 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_9_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_0_109 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_22_3 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_14_29 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_6_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_17 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_28 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_39 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
Xoutput3 net3 vss vss vcc vcc reg_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_22_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_22_29 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XANTENNA_input1_A spi_mosi vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_10_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_69_ clknet_1_1__leaf_spi_clk _03_ _13_ vss vss vcc vcc t\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_23_61 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_0_21 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_15_3 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_20_62 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_20_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_6_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_18 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_29 vss vss vcc vcc sky130_fd_sc_hd__decap_3
Xoutput4 net4 vss vss vcc vcc reg_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_14_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_68_ clknet_1_1__leaf_spi_clk _02_ _12_ vss vss vcc vcc t\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_2_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_62 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_19 vss vss vcc vcc sky130_fd_sc_hd__decap_3
Xoutput5 net5 vss vss vcc vcc reg_addr[2] sky130_fd_sc_hd__buf_2
XTAP_110 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_22_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_9_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_12_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_67_ _01_ _11_ vss vss vcc vcc net5 sky130_fd_sc_hd__dlxtn_1
XFILLER_5_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_2_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_74 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_18_41 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_20_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_6_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
Xoutput6 net6 vss vss vcc vcc reg_clk sky130_fd_sc_hd__buf_2
XFILLER_15_20 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XTAP_111 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
.ends

