magic
tech sky130B
magscale 1 2
timestamp 1675783699
<< viali >>
rect 1869 21641 1903 21675
rect 4813 21641 4847 21675
rect 7757 21641 7791 21675
rect 10701 21641 10735 21675
rect 14381 21641 14415 21675
rect 16957 21641 16991 21675
rect 19533 21641 19567 21675
rect 22201 21641 22235 21675
rect 2053 21505 2087 21539
rect 4997 21505 5031 21539
rect 7941 21505 7975 21539
rect 10885 21505 10919 21539
rect 14565 21505 14599 21539
rect 17141 21505 17175 21539
rect 19717 21505 19751 21539
rect 22017 21505 22051 21539
rect 2513 21301 2547 21335
rect 5549 21301 5583 21335
rect 8401 21301 8435 21335
rect 11713 21301 11747 21335
rect 17877 14025 17911 14059
rect 17141 13889 17175 13923
rect 16865 13821 16899 13855
rect 16681 13277 16715 13311
rect 16957 13277 16991 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 17693 13141 17727 13175
rect 18705 13141 18739 13175
rect 16221 12937 16255 12971
rect 16865 12937 16899 12971
rect 16129 12801 16163 12835
rect 16313 12801 16347 12835
rect 16865 12801 16899 12835
rect 17049 12801 17083 12835
rect 18797 12801 18831 12835
rect 19073 12801 19107 12835
rect 19809 12801 19843 12835
rect 19993 12801 20027 12835
rect 18935 12733 18969 12767
rect 19349 12665 19383 12699
rect 18153 12597 18187 12631
rect 18429 12393 18463 12427
rect 20453 12393 20487 12427
rect 18613 12325 18647 12359
rect 15577 12257 15611 12291
rect 16129 12257 16163 12291
rect 19441 12257 19475 12291
rect 15485 12189 15519 12223
rect 15669 12189 15703 12223
rect 16405 12189 16439 12223
rect 19717 12189 19751 12223
rect 18889 12121 18923 12155
rect 17141 12053 17175 12087
rect 17969 11849 18003 11883
rect 17233 11713 17267 11747
rect 16957 11645 16991 11679
rect 18889 11645 18923 11679
rect 18613 11577 18647 11611
rect 18429 11509 18463 11543
rect 17233 11305 17267 11339
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 17785 11101 17819 11135
rect 17969 11101 18003 11135
rect 17877 10965 17911 10999
rect 17601 10625 17635 10659
rect 17877 10625 17911 10659
rect 18889 10625 18923 10659
rect 21189 10625 21223 10659
rect 18613 10557 18647 10591
rect 21005 10557 21039 10591
rect 16865 10421 16899 10455
rect 19625 10421 19659 10455
rect 20085 10421 20119 10455
rect 21373 10421 21407 10455
rect 20453 10217 20487 10251
rect 17693 10149 17727 10183
rect 17233 10081 17267 10115
rect 17969 10081 18003 10115
rect 18086 10081 18120 10115
rect 18245 10081 18279 10115
rect 21281 10081 21315 10115
rect 21557 10081 21591 10115
rect 17049 10013 17083 10047
rect 19441 10013 19475 10047
rect 19717 10013 19751 10047
rect 16589 9877 16623 9911
rect 18889 9877 18923 9911
rect 18153 9673 18187 9707
rect 18797 9673 18831 9707
rect 19441 9673 19475 9707
rect 19993 9673 20027 9707
rect 18705 9537 18739 9571
rect 18889 9537 18923 9571
rect 19349 9537 19383 9571
rect 19533 9537 19567 9571
rect 21005 9537 21039 9571
rect 21189 9537 21223 9571
rect 21097 9469 21131 9503
rect 22017 8517 22051 8551
rect 19165 8449 19199 8483
rect 20269 8449 20303 8483
rect 21189 8449 21223 8483
rect 22201 8449 22235 8483
rect 22293 8449 22327 8483
rect 20545 8381 20579 8415
rect 21465 8381 21499 8415
rect 18705 8313 18739 8347
rect 20361 8313 20395 8347
rect 21005 8313 21039 8347
rect 22017 8313 22051 8347
rect 18889 8245 18923 8279
rect 20453 8245 20487 8279
rect 21373 8245 21407 8279
rect 18061 7837 18095 7871
rect 18429 7837 18463 7871
rect 18889 7837 18923 7871
rect 19441 7837 19475 7871
rect 18613 7769 18647 7803
rect 19625 7769 19659 7803
rect 19809 7701 19843 7735
rect 18797 7497 18831 7531
rect 18613 7361 18647 7395
rect 18889 7361 18923 7395
rect 18429 7293 18463 7327
rect 21465 6409 21499 6443
rect 20352 6341 20386 6375
rect 20085 6205 20119 6239
rect 20085 5661 20119 5695
rect 20330 5593 20364 5627
rect 21465 5525 21499 5559
rect 20637 5321 20671 5355
rect 19993 5253 20027 5287
rect 20545 5185 20579 5219
rect 18705 4981 18739 5015
rect 18889 4777 18923 4811
rect 20269 4777 20303 4811
rect 18245 4641 18279 4675
rect 18403 4573 18437 4607
rect 18613 4573 18647 4607
rect 18705 4573 18739 4607
rect 19441 4573 19475 4607
rect 19625 4573 19659 4607
rect 21649 4573 21683 4607
rect 18521 4505 18555 4539
rect 19533 4505 19567 4539
rect 21404 4505 21438 4539
rect 22201 4437 22235 4471
rect 19349 4097 19383 4131
rect 20249 4097 20283 4131
rect 22017 4097 22051 4131
rect 19441 4029 19475 4063
rect 19993 4029 20027 4063
rect 21373 3893 21407 3927
rect 18337 3689 18371 3723
rect 20821 3689 20855 3723
rect 18153 3485 18187 3519
rect 18337 3485 18371 3519
rect 22293 3417 22327 3451
rect 13185 3145 13219 3179
rect 22109 3145 22143 3179
rect 13001 3009 13035 3043
rect 13369 3009 13403 3043
rect 13645 3009 13679 3043
rect 14105 3009 14139 3043
rect 14381 3009 14415 3043
rect 15577 3009 15611 3043
rect 16865 3009 16899 3043
rect 17877 3009 17911 3043
rect 22017 3009 22051 3043
rect 14197 2941 14231 2975
rect 18061 2941 18095 2975
rect 18337 2941 18371 2975
rect 14565 2873 14599 2907
rect 15761 2873 15795 2907
rect 17049 2873 17083 2907
rect 13461 2805 13495 2839
rect 14289 2805 14323 2839
rect 10241 2601 10275 2635
rect 14289 2601 14323 2635
rect 17509 2601 17543 2635
rect 2329 2533 2363 2567
rect 18889 2465 18923 2499
rect 22109 2465 22143 2499
rect 2145 2397 2179 2431
rect 2789 2397 2823 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 19717 2397 19751 2431
rect 21465 2397 21499 2431
rect 22017 2397 22051 2431
rect 18644 2329 18678 2363
rect 6745 2261 6779 2295
<< metal1 >>
rect 1104 21786 22976 21808
rect 1104 21734 6378 21786
rect 6430 21734 6442 21786
rect 6494 21734 6506 21786
rect 6558 21734 6570 21786
rect 6622 21734 6634 21786
rect 6686 21734 11806 21786
rect 11858 21734 11870 21786
rect 11922 21734 11934 21786
rect 11986 21734 11998 21786
rect 12050 21734 12062 21786
rect 12114 21734 17234 21786
rect 17286 21734 17298 21786
rect 17350 21734 17362 21786
rect 17414 21734 17426 21786
rect 17478 21734 17490 21786
rect 17542 21734 22662 21786
rect 22714 21734 22726 21786
rect 22778 21734 22790 21786
rect 22842 21734 22854 21786
rect 22906 21734 22918 21786
rect 22970 21734 22976 21786
rect 1104 21712 22976 21734
rect 1854 21672 1860 21684
rect 1815 21644 1860 21672
rect 1854 21632 1860 21644
rect 1912 21632 1918 21684
rect 4798 21672 4804 21684
rect 4759 21644 4804 21672
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 7742 21672 7748 21684
rect 7703 21644 7748 21672
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 10686 21672 10692 21684
rect 10647 21644 10692 21672
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 13814 21632 13820 21684
rect 13872 21672 13878 21684
rect 14369 21675 14427 21681
rect 14369 21672 14381 21675
rect 13872 21644 14381 21672
rect 13872 21632 13878 21644
rect 14369 21641 14381 21644
rect 14415 21641 14427 21675
rect 14369 21635 14427 21641
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 16945 21675 17003 21681
rect 16945 21672 16957 21675
rect 16632 21644 16957 21672
rect 16632 21632 16638 21644
rect 16945 21641 16957 21644
rect 16991 21641 17003 21675
rect 19518 21672 19524 21684
rect 19479 21644 19524 21672
rect 16945 21635 17003 21641
rect 19518 21632 19524 21644
rect 19576 21632 19582 21684
rect 22186 21672 22192 21684
rect 22147 21644 22192 21672
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21536 2099 21539
rect 2498 21536 2504 21548
rect 2087 21508 2504 21536
rect 2087 21505 2099 21508
rect 2041 21499 2099 21505
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21536 5043 21539
rect 7929 21539 7987 21545
rect 5031 21508 5580 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 2498 21332 2504 21344
rect 2459 21304 2504 21332
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 5552 21341 5580 21508
rect 7929 21505 7941 21539
rect 7975 21536 7987 21539
rect 8386 21536 8392 21548
rect 7975 21508 8392 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 8386 21496 8392 21508
rect 8444 21496 8450 21548
rect 10873 21539 10931 21545
rect 10873 21505 10885 21539
rect 10919 21536 10931 21539
rect 11698 21536 11704 21548
rect 10919 21508 11704 21536
rect 10919 21505 10931 21508
rect 10873 21499 10931 21505
rect 11698 21496 11704 21508
rect 11756 21496 11762 21548
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 17129 21539 17187 21545
rect 14599 21508 16574 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 16546 21468 16574 21508
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 17862 21536 17868 21548
rect 17175 21508 17868 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21536 19763 21539
rect 20438 21536 20444 21548
rect 19751 21508 20444 21536
rect 19751 21505 19763 21508
rect 19705 21499 19763 21505
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 19058 21468 19064 21480
rect 16546 21440 19064 21468
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 19794 21428 19800 21480
rect 19852 21468 19858 21480
rect 22020 21468 22048 21499
rect 19852 21440 22048 21468
rect 19852 21428 19858 21440
rect 5537 21335 5595 21341
rect 5537 21301 5549 21335
rect 5583 21332 5595 21335
rect 6178 21332 6184 21344
rect 5583 21304 6184 21332
rect 5583 21301 5595 21304
rect 5537 21295 5595 21301
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 8386 21332 8392 21344
rect 8347 21304 8392 21332
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 11698 21332 11704 21344
rect 11659 21304 11704 21332
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 1104 21242 22816 21264
rect 1104 21190 3664 21242
rect 3716 21190 3728 21242
rect 3780 21190 3792 21242
rect 3844 21190 3856 21242
rect 3908 21190 3920 21242
rect 3972 21190 9092 21242
rect 9144 21190 9156 21242
rect 9208 21190 9220 21242
rect 9272 21190 9284 21242
rect 9336 21190 9348 21242
rect 9400 21190 14520 21242
rect 14572 21190 14584 21242
rect 14636 21190 14648 21242
rect 14700 21190 14712 21242
rect 14764 21190 14776 21242
rect 14828 21190 19948 21242
rect 20000 21190 20012 21242
rect 20064 21190 20076 21242
rect 20128 21190 20140 21242
rect 20192 21190 20204 21242
rect 20256 21190 22816 21242
rect 1104 21168 22816 21190
rect 1104 20698 22976 20720
rect 1104 20646 6378 20698
rect 6430 20646 6442 20698
rect 6494 20646 6506 20698
rect 6558 20646 6570 20698
rect 6622 20646 6634 20698
rect 6686 20646 11806 20698
rect 11858 20646 11870 20698
rect 11922 20646 11934 20698
rect 11986 20646 11998 20698
rect 12050 20646 12062 20698
rect 12114 20646 17234 20698
rect 17286 20646 17298 20698
rect 17350 20646 17362 20698
rect 17414 20646 17426 20698
rect 17478 20646 17490 20698
rect 17542 20646 22662 20698
rect 22714 20646 22726 20698
rect 22778 20646 22790 20698
rect 22842 20646 22854 20698
rect 22906 20646 22918 20698
rect 22970 20646 22976 20698
rect 1104 20624 22976 20646
rect 1104 20154 22816 20176
rect 1104 20102 3664 20154
rect 3716 20102 3728 20154
rect 3780 20102 3792 20154
rect 3844 20102 3856 20154
rect 3908 20102 3920 20154
rect 3972 20102 9092 20154
rect 9144 20102 9156 20154
rect 9208 20102 9220 20154
rect 9272 20102 9284 20154
rect 9336 20102 9348 20154
rect 9400 20102 14520 20154
rect 14572 20102 14584 20154
rect 14636 20102 14648 20154
rect 14700 20102 14712 20154
rect 14764 20102 14776 20154
rect 14828 20102 19948 20154
rect 20000 20102 20012 20154
rect 20064 20102 20076 20154
rect 20128 20102 20140 20154
rect 20192 20102 20204 20154
rect 20256 20102 22816 20154
rect 1104 20080 22816 20102
rect 1104 19610 22976 19632
rect 1104 19558 6378 19610
rect 6430 19558 6442 19610
rect 6494 19558 6506 19610
rect 6558 19558 6570 19610
rect 6622 19558 6634 19610
rect 6686 19558 11806 19610
rect 11858 19558 11870 19610
rect 11922 19558 11934 19610
rect 11986 19558 11998 19610
rect 12050 19558 12062 19610
rect 12114 19558 17234 19610
rect 17286 19558 17298 19610
rect 17350 19558 17362 19610
rect 17414 19558 17426 19610
rect 17478 19558 17490 19610
rect 17542 19558 22662 19610
rect 22714 19558 22726 19610
rect 22778 19558 22790 19610
rect 22842 19558 22854 19610
rect 22906 19558 22918 19610
rect 22970 19558 22976 19610
rect 1104 19536 22976 19558
rect 1104 19066 22816 19088
rect 1104 19014 3664 19066
rect 3716 19014 3728 19066
rect 3780 19014 3792 19066
rect 3844 19014 3856 19066
rect 3908 19014 3920 19066
rect 3972 19014 9092 19066
rect 9144 19014 9156 19066
rect 9208 19014 9220 19066
rect 9272 19014 9284 19066
rect 9336 19014 9348 19066
rect 9400 19014 14520 19066
rect 14572 19014 14584 19066
rect 14636 19014 14648 19066
rect 14700 19014 14712 19066
rect 14764 19014 14776 19066
rect 14828 19014 19948 19066
rect 20000 19014 20012 19066
rect 20064 19014 20076 19066
rect 20128 19014 20140 19066
rect 20192 19014 20204 19066
rect 20256 19014 22816 19066
rect 1104 18992 22816 19014
rect 1104 18522 22976 18544
rect 1104 18470 6378 18522
rect 6430 18470 6442 18522
rect 6494 18470 6506 18522
rect 6558 18470 6570 18522
rect 6622 18470 6634 18522
rect 6686 18470 11806 18522
rect 11858 18470 11870 18522
rect 11922 18470 11934 18522
rect 11986 18470 11998 18522
rect 12050 18470 12062 18522
rect 12114 18470 17234 18522
rect 17286 18470 17298 18522
rect 17350 18470 17362 18522
rect 17414 18470 17426 18522
rect 17478 18470 17490 18522
rect 17542 18470 22662 18522
rect 22714 18470 22726 18522
rect 22778 18470 22790 18522
rect 22842 18470 22854 18522
rect 22906 18470 22918 18522
rect 22970 18470 22976 18522
rect 1104 18448 22976 18470
rect 1104 17978 22816 18000
rect 1104 17926 3664 17978
rect 3716 17926 3728 17978
rect 3780 17926 3792 17978
rect 3844 17926 3856 17978
rect 3908 17926 3920 17978
rect 3972 17926 9092 17978
rect 9144 17926 9156 17978
rect 9208 17926 9220 17978
rect 9272 17926 9284 17978
rect 9336 17926 9348 17978
rect 9400 17926 14520 17978
rect 14572 17926 14584 17978
rect 14636 17926 14648 17978
rect 14700 17926 14712 17978
rect 14764 17926 14776 17978
rect 14828 17926 19948 17978
rect 20000 17926 20012 17978
rect 20064 17926 20076 17978
rect 20128 17926 20140 17978
rect 20192 17926 20204 17978
rect 20256 17926 22816 17978
rect 1104 17904 22816 17926
rect 1104 17434 22976 17456
rect 1104 17382 6378 17434
rect 6430 17382 6442 17434
rect 6494 17382 6506 17434
rect 6558 17382 6570 17434
rect 6622 17382 6634 17434
rect 6686 17382 11806 17434
rect 11858 17382 11870 17434
rect 11922 17382 11934 17434
rect 11986 17382 11998 17434
rect 12050 17382 12062 17434
rect 12114 17382 17234 17434
rect 17286 17382 17298 17434
rect 17350 17382 17362 17434
rect 17414 17382 17426 17434
rect 17478 17382 17490 17434
rect 17542 17382 22662 17434
rect 22714 17382 22726 17434
rect 22778 17382 22790 17434
rect 22842 17382 22854 17434
rect 22906 17382 22918 17434
rect 22970 17382 22976 17434
rect 1104 17360 22976 17382
rect 1104 16890 22816 16912
rect 1104 16838 3664 16890
rect 3716 16838 3728 16890
rect 3780 16838 3792 16890
rect 3844 16838 3856 16890
rect 3908 16838 3920 16890
rect 3972 16838 9092 16890
rect 9144 16838 9156 16890
rect 9208 16838 9220 16890
rect 9272 16838 9284 16890
rect 9336 16838 9348 16890
rect 9400 16838 14520 16890
rect 14572 16838 14584 16890
rect 14636 16838 14648 16890
rect 14700 16838 14712 16890
rect 14764 16838 14776 16890
rect 14828 16838 19948 16890
rect 20000 16838 20012 16890
rect 20064 16838 20076 16890
rect 20128 16838 20140 16890
rect 20192 16838 20204 16890
rect 20256 16838 22816 16890
rect 1104 16816 22816 16838
rect 1104 16346 22976 16368
rect 1104 16294 6378 16346
rect 6430 16294 6442 16346
rect 6494 16294 6506 16346
rect 6558 16294 6570 16346
rect 6622 16294 6634 16346
rect 6686 16294 11806 16346
rect 11858 16294 11870 16346
rect 11922 16294 11934 16346
rect 11986 16294 11998 16346
rect 12050 16294 12062 16346
rect 12114 16294 17234 16346
rect 17286 16294 17298 16346
rect 17350 16294 17362 16346
rect 17414 16294 17426 16346
rect 17478 16294 17490 16346
rect 17542 16294 22662 16346
rect 22714 16294 22726 16346
rect 22778 16294 22790 16346
rect 22842 16294 22854 16346
rect 22906 16294 22918 16346
rect 22970 16294 22976 16346
rect 1104 16272 22976 16294
rect 1104 15802 22816 15824
rect 1104 15750 3664 15802
rect 3716 15750 3728 15802
rect 3780 15750 3792 15802
rect 3844 15750 3856 15802
rect 3908 15750 3920 15802
rect 3972 15750 9092 15802
rect 9144 15750 9156 15802
rect 9208 15750 9220 15802
rect 9272 15750 9284 15802
rect 9336 15750 9348 15802
rect 9400 15750 14520 15802
rect 14572 15750 14584 15802
rect 14636 15750 14648 15802
rect 14700 15750 14712 15802
rect 14764 15750 14776 15802
rect 14828 15750 19948 15802
rect 20000 15750 20012 15802
rect 20064 15750 20076 15802
rect 20128 15750 20140 15802
rect 20192 15750 20204 15802
rect 20256 15750 22816 15802
rect 1104 15728 22816 15750
rect 1104 15258 22976 15280
rect 1104 15206 6378 15258
rect 6430 15206 6442 15258
rect 6494 15206 6506 15258
rect 6558 15206 6570 15258
rect 6622 15206 6634 15258
rect 6686 15206 11806 15258
rect 11858 15206 11870 15258
rect 11922 15206 11934 15258
rect 11986 15206 11998 15258
rect 12050 15206 12062 15258
rect 12114 15206 17234 15258
rect 17286 15206 17298 15258
rect 17350 15206 17362 15258
rect 17414 15206 17426 15258
rect 17478 15206 17490 15258
rect 17542 15206 22662 15258
rect 22714 15206 22726 15258
rect 22778 15206 22790 15258
rect 22842 15206 22854 15258
rect 22906 15206 22918 15258
rect 22970 15206 22976 15258
rect 1104 15184 22976 15206
rect 1104 14714 22816 14736
rect 1104 14662 3664 14714
rect 3716 14662 3728 14714
rect 3780 14662 3792 14714
rect 3844 14662 3856 14714
rect 3908 14662 3920 14714
rect 3972 14662 9092 14714
rect 9144 14662 9156 14714
rect 9208 14662 9220 14714
rect 9272 14662 9284 14714
rect 9336 14662 9348 14714
rect 9400 14662 14520 14714
rect 14572 14662 14584 14714
rect 14636 14662 14648 14714
rect 14700 14662 14712 14714
rect 14764 14662 14776 14714
rect 14828 14662 19948 14714
rect 20000 14662 20012 14714
rect 20064 14662 20076 14714
rect 20128 14662 20140 14714
rect 20192 14662 20204 14714
rect 20256 14662 22816 14714
rect 1104 14640 22816 14662
rect 1104 14170 22976 14192
rect 1104 14118 6378 14170
rect 6430 14118 6442 14170
rect 6494 14118 6506 14170
rect 6558 14118 6570 14170
rect 6622 14118 6634 14170
rect 6686 14118 11806 14170
rect 11858 14118 11870 14170
rect 11922 14118 11934 14170
rect 11986 14118 11998 14170
rect 12050 14118 12062 14170
rect 12114 14118 17234 14170
rect 17286 14118 17298 14170
rect 17350 14118 17362 14170
rect 17414 14118 17426 14170
rect 17478 14118 17490 14170
rect 17542 14118 22662 14170
rect 22714 14118 22726 14170
rect 22778 14118 22790 14170
rect 22842 14118 22854 14170
rect 22906 14118 22918 14170
rect 22970 14118 22976 14170
rect 1104 14096 22976 14118
rect 17862 14056 17868 14068
rect 17823 14028 17868 14056
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17129 13923 17187 13929
rect 17129 13920 17141 13923
rect 17092 13892 17141 13920
rect 17092 13880 17098 13892
rect 17129 13889 17141 13892
rect 17175 13889 17187 13923
rect 17129 13883 17187 13889
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 1104 13626 22816 13648
rect 1104 13574 3664 13626
rect 3716 13574 3728 13626
rect 3780 13574 3792 13626
rect 3844 13574 3856 13626
rect 3908 13574 3920 13626
rect 3972 13574 9092 13626
rect 9144 13574 9156 13626
rect 9208 13574 9220 13626
rect 9272 13574 9284 13626
rect 9336 13574 9348 13626
rect 9400 13574 14520 13626
rect 14572 13574 14584 13626
rect 14636 13574 14648 13626
rect 14700 13574 14712 13626
rect 14764 13574 14776 13626
rect 14828 13574 19948 13626
rect 20000 13574 20012 13626
rect 20064 13574 20076 13626
rect 20128 13574 20140 13626
rect 20192 13574 20204 13626
rect 20256 13574 22816 13626
rect 1104 13552 22816 13574
rect 16206 13268 16212 13320
rect 16264 13308 16270 13320
rect 16669 13311 16727 13317
rect 16669 13308 16681 13311
rect 16264 13280 16681 13308
rect 16264 13268 16270 13280
rect 16669 13277 16681 13280
rect 16715 13277 16727 13311
rect 16942 13308 16948 13320
rect 16903 13280 16948 13308
rect 16669 13271 16727 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18509 13311 18567 13317
rect 18509 13308 18521 13311
rect 18012 13280 18521 13308
rect 18012 13268 18018 13280
rect 18509 13277 18521 13280
rect 18555 13277 18567 13311
rect 18690 13308 18696 13320
rect 18651 13280 18696 13308
rect 18509 13271 18567 13277
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 17678 13172 17684 13184
rect 8444 13144 17684 13172
rect 8444 13132 8450 13144
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 18693 13175 18751 13181
rect 18693 13141 18705 13175
rect 18739 13172 18751 13175
rect 19426 13172 19432 13184
rect 18739 13144 19432 13172
rect 18739 13141 18751 13144
rect 18693 13135 18751 13141
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 1104 13082 22976 13104
rect 1104 13030 6378 13082
rect 6430 13030 6442 13082
rect 6494 13030 6506 13082
rect 6558 13030 6570 13082
rect 6622 13030 6634 13082
rect 6686 13030 11806 13082
rect 11858 13030 11870 13082
rect 11922 13030 11934 13082
rect 11986 13030 11998 13082
rect 12050 13030 12062 13082
rect 12114 13030 17234 13082
rect 17286 13030 17298 13082
rect 17350 13030 17362 13082
rect 17414 13030 17426 13082
rect 17478 13030 17490 13082
rect 17542 13030 22662 13082
rect 22714 13030 22726 13082
rect 22778 13030 22790 13082
rect 22842 13030 22854 13082
rect 22906 13030 22918 13082
rect 22970 13030 22976 13082
rect 1104 13008 22976 13030
rect 16206 12968 16212 12980
rect 16167 12940 16212 12968
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 16114 12832 16120 12844
rect 16075 12804 16120 12832
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16850 12832 16856 12844
rect 16347 12804 16574 12832
rect 16811 12804 16856 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16546 12696 16574 12804
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17954 12832 17960 12844
rect 17083 12804 17960 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 18782 12792 18788 12844
rect 18840 12832 18846 12844
rect 19058 12832 19064 12844
rect 18840 12804 18885 12832
rect 19019 12804 19064 12832
rect 18840 12792 18846 12804
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 19794 12832 19800 12844
rect 19755 12804 19800 12832
rect 19794 12792 19800 12804
rect 19852 12792 19858 12844
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12832 20039 12835
rect 20438 12832 20444 12844
rect 20027 12804 20444 12832
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 18923 12767 18981 12773
rect 18923 12764 18935 12767
rect 17920 12736 18935 12764
rect 17920 12724 17926 12736
rect 18923 12733 18935 12736
rect 18969 12733 18981 12767
rect 18923 12727 18981 12733
rect 19337 12699 19395 12705
rect 16546 12668 18276 12696
rect 18138 12628 18144 12640
rect 18099 12600 18144 12628
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 18248 12628 18276 12668
rect 19337 12665 19349 12699
rect 19383 12665 19395 12699
rect 19337 12659 19395 12665
rect 18690 12628 18696 12640
rect 18248 12600 18696 12628
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 18966 12588 18972 12640
rect 19024 12628 19030 12640
rect 19352 12628 19380 12659
rect 19024 12600 19380 12628
rect 19024 12588 19030 12600
rect 1104 12538 22816 12560
rect 1104 12486 3664 12538
rect 3716 12486 3728 12538
rect 3780 12486 3792 12538
rect 3844 12486 3856 12538
rect 3908 12486 3920 12538
rect 3972 12486 9092 12538
rect 9144 12486 9156 12538
rect 9208 12486 9220 12538
rect 9272 12486 9284 12538
rect 9336 12486 9348 12538
rect 9400 12486 14520 12538
rect 14572 12486 14584 12538
rect 14636 12486 14648 12538
rect 14700 12486 14712 12538
rect 14764 12486 14776 12538
rect 14828 12486 19948 12538
rect 20000 12486 20012 12538
rect 20064 12486 20076 12538
rect 20128 12486 20140 12538
rect 20192 12486 20204 12538
rect 20256 12486 22816 12538
rect 1104 12464 22816 12486
rect 16114 12384 16120 12436
rect 16172 12424 16178 12436
rect 18230 12424 18236 12436
rect 16172 12396 18236 12424
rect 16172 12384 16178 12396
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 18417 12427 18475 12433
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 18690 12424 18696 12436
rect 18463 12396 18696 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 20438 12424 20444 12436
rect 20399 12396 20444 12424
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 18601 12359 18659 12365
rect 18601 12325 18613 12359
rect 18647 12356 18659 12359
rect 18874 12356 18880 12368
rect 18647 12328 18880 12356
rect 18647 12325 18659 12328
rect 18601 12319 18659 12325
rect 18874 12316 18880 12328
rect 18932 12316 18938 12368
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12288 15623 12291
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 15611 12260 16129 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 19426 12288 19432 12300
rect 19387 12260 19432 12288
rect 16117 12251 16175 12257
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12189 15531 12223
rect 15473 12183 15531 12189
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 16022 12220 16028 12232
rect 15703 12192 16028 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 15488 12152 15516 12183
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16942 12220 16948 12232
rect 16439 12192 16948 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 19702 12220 19708 12232
rect 19663 12192 19708 12220
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 16850 12152 16856 12164
rect 15488 12124 16856 12152
rect 16850 12112 16856 12124
rect 16908 12112 16914 12164
rect 18782 12112 18788 12164
rect 18840 12152 18846 12164
rect 18877 12155 18935 12161
rect 18877 12152 18889 12155
rect 18840 12124 18889 12152
rect 18840 12112 18846 12124
rect 18877 12121 18889 12124
rect 18923 12152 18935 12155
rect 18966 12152 18972 12164
rect 18923 12124 18972 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 18966 12112 18972 12124
rect 19024 12112 19030 12164
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 17129 12087 17187 12093
rect 17129 12084 17141 12087
rect 6236 12056 17141 12084
rect 6236 12044 6242 12056
rect 17129 12053 17141 12056
rect 17175 12084 17187 12087
rect 18046 12084 18052 12096
rect 17175 12056 18052 12084
rect 17175 12053 17187 12056
rect 17129 12047 17187 12053
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 1104 11994 22976 12016
rect 1104 11942 6378 11994
rect 6430 11942 6442 11994
rect 6494 11942 6506 11994
rect 6558 11942 6570 11994
rect 6622 11942 6634 11994
rect 6686 11942 11806 11994
rect 11858 11942 11870 11994
rect 11922 11942 11934 11994
rect 11986 11942 11998 11994
rect 12050 11942 12062 11994
rect 12114 11942 17234 11994
rect 17286 11942 17298 11994
rect 17350 11942 17362 11994
rect 17414 11942 17426 11994
rect 17478 11942 17490 11994
rect 17542 11942 22662 11994
rect 22714 11942 22726 11994
rect 22778 11942 22790 11994
rect 22842 11942 22854 11994
rect 22906 11942 22918 11994
rect 22970 11942 22976 11994
rect 1104 11920 22976 11942
rect 17957 11883 18015 11889
rect 17957 11849 17969 11883
rect 18003 11880 18015 11883
rect 19058 11880 19064 11892
rect 18003 11852 19064 11880
rect 18003 11849 18015 11852
rect 17957 11843 18015 11849
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 16942 11772 16948 11824
rect 17000 11772 17006 11824
rect 16960 11744 16988 11772
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16960 11716 17233 11744
rect 17221 11713 17233 11716
rect 17267 11744 17279 11747
rect 17586 11744 17592 11756
rect 17267 11716 17592 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 16942 11676 16948 11688
rect 16903 11648 16948 11676
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 18874 11676 18880 11688
rect 18835 11648 18880 11676
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 18601 11611 18659 11617
rect 18601 11577 18613 11611
rect 18647 11608 18659 11611
rect 18966 11608 18972 11620
rect 18647 11580 18972 11608
rect 18647 11577 18659 11580
rect 18601 11571 18659 11577
rect 18966 11568 18972 11580
rect 19024 11568 19030 11620
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 18417 11543 18475 11549
rect 18417 11540 18429 11543
rect 16908 11512 18429 11540
rect 16908 11500 16914 11512
rect 18417 11509 18429 11512
rect 18463 11509 18475 11543
rect 18417 11503 18475 11509
rect 1104 11450 22816 11472
rect 1104 11398 3664 11450
rect 3716 11398 3728 11450
rect 3780 11398 3792 11450
rect 3844 11398 3856 11450
rect 3908 11398 3920 11450
rect 3972 11398 9092 11450
rect 9144 11398 9156 11450
rect 9208 11398 9220 11450
rect 9272 11398 9284 11450
rect 9336 11398 9348 11450
rect 9400 11398 14520 11450
rect 14572 11398 14584 11450
rect 14636 11398 14648 11450
rect 14700 11398 14712 11450
rect 14764 11398 14776 11450
rect 14828 11398 19948 11450
rect 20000 11398 20012 11450
rect 20064 11398 20076 11450
rect 20128 11398 20140 11450
rect 20192 11398 20204 11450
rect 20256 11398 22816 11450
rect 1104 11376 22816 11398
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 17000 11308 17233 11336
rect 17000 11296 17006 11308
rect 17221 11305 17233 11308
rect 17267 11305 17279 11339
rect 17221 11299 17279 11305
rect 21542 11268 21548 11280
rect 17696 11240 21548 11268
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11132 17371 11135
rect 17696 11132 17724 11240
rect 21542 11228 21548 11240
rect 21600 11228 21606 11280
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 17359 11104 17785 11132
rect 17359 11101 17371 11104
rect 17313 11095 17371 11101
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 18230 11132 18236 11144
rect 18003 11104 18236 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 17144 11064 17172 11095
rect 18230 11092 18236 11104
rect 18288 11132 18294 11144
rect 18690 11132 18696 11144
rect 18288 11104 18696 11132
rect 18288 11092 18294 11104
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 19242 11064 19248 11076
rect 17144 11036 19248 11064
rect 17972 11008 18000 11036
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 17862 10996 17868 11008
rect 17823 10968 17868 10996
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 17954 10956 17960 11008
rect 18012 10956 18018 11008
rect 1104 10906 22976 10928
rect 1104 10854 6378 10906
rect 6430 10854 6442 10906
rect 6494 10854 6506 10906
rect 6558 10854 6570 10906
rect 6622 10854 6634 10906
rect 6686 10854 11806 10906
rect 11858 10854 11870 10906
rect 11922 10854 11934 10906
rect 11986 10854 11998 10906
rect 12050 10854 12062 10906
rect 12114 10854 17234 10906
rect 17286 10854 17298 10906
rect 17350 10854 17362 10906
rect 17414 10854 17426 10906
rect 17478 10854 17490 10906
rect 17542 10854 22662 10906
rect 22714 10854 22726 10906
rect 22778 10854 22790 10906
rect 22842 10854 22854 10906
rect 22906 10854 22918 10906
rect 22970 10854 22976 10906
rect 1104 10832 22976 10854
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 18932 10764 21220 10792
rect 18932 10752 18938 10764
rect 19702 10724 19708 10736
rect 17696 10696 19708 10724
rect 17586 10656 17592 10668
rect 17499 10628 17592 10656
rect 17586 10616 17592 10628
rect 17644 10656 17650 10668
rect 17696 10656 17724 10696
rect 17862 10656 17868 10668
rect 17644 10628 17724 10656
rect 17823 10628 17868 10656
rect 17644 10616 17650 10628
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 18892 10665 18920 10696
rect 19702 10684 19708 10696
rect 19760 10684 19766 10736
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 18966 10616 18972 10668
rect 19024 10656 19030 10668
rect 21192 10665 21220 10764
rect 21177 10659 21235 10665
rect 19024 10628 21036 10656
rect 19024 10616 19030 10628
rect 18598 10588 18604 10600
rect 18559 10560 18604 10588
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 21008 10597 21036 10628
rect 21177 10625 21189 10659
rect 21223 10656 21235 10659
rect 21358 10656 21364 10668
rect 21223 10628 21364 10656
rect 21223 10625 21235 10628
rect 21177 10619 21235 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10557 21051 10591
rect 20993 10551 21051 10557
rect 21008 10520 21036 10551
rect 21174 10520 21180 10532
rect 21008 10492 21180 10520
rect 21174 10480 21180 10492
rect 21232 10480 21238 10532
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 17276 10424 19625 10452
rect 17276 10412 17282 10424
rect 19613 10421 19625 10424
rect 19659 10452 19671 10455
rect 20073 10455 20131 10461
rect 20073 10452 20085 10455
rect 19659 10424 20085 10452
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 20073 10421 20085 10424
rect 20119 10421 20131 10455
rect 20073 10415 20131 10421
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21361 10455 21419 10461
rect 21361 10452 21373 10455
rect 21324 10424 21373 10452
rect 21324 10412 21330 10424
rect 21361 10421 21373 10424
rect 21407 10421 21419 10455
rect 21361 10415 21419 10421
rect 1104 10362 22816 10384
rect 1104 10310 3664 10362
rect 3716 10310 3728 10362
rect 3780 10310 3792 10362
rect 3844 10310 3856 10362
rect 3908 10310 3920 10362
rect 3972 10310 9092 10362
rect 9144 10310 9156 10362
rect 9208 10310 9220 10362
rect 9272 10310 9284 10362
rect 9336 10310 9348 10362
rect 9400 10310 14520 10362
rect 14572 10310 14584 10362
rect 14636 10310 14648 10362
rect 14700 10310 14712 10362
rect 14764 10310 14776 10362
rect 14828 10310 19948 10362
rect 20000 10310 20012 10362
rect 20064 10310 20076 10362
rect 20128 10310 20140 10362
rect 20192 10310 20204 10362
rect 20256 10310 22816 10362
rect 1104 10288 22816 10310
rect 18874 10248 18880 10260
rect 17788 10220 18880 10248
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 17681 10183 17739 10189
rect 16908 10152 17356 10180
rect 16908 10140 16914 10152
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 17218 10112 17224 10124
rect 11756 10084 17224 10112
rect 11756 10072 11762 10084
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17328 10112 17356 10152
rect 17681 10149 17693 10183
rect 17727 10180 17739 10183
rect 17788 10180 17816 10220
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 19794 10208 19800 10260
rect 19852 10248 19858 10260
rect 20441 10251 20499 10257
rect 20441 10248 20453 10251
rect 19852 10220 20453 10248
rect 19852 10208 19858 10220
rect 20441 10217 20453 10220
rect 20487 10217 20499 10251
rect 20441 10211 20499 10217
rect 17727 10152 17816 10180
rect 17727 10149 17739 10152
rect 17681 10143 17739 10149
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 17328 10084 17969 10112
rect 17957 10081 17969 10084
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 18046 10072 18052 10124
rect 18104 10121 18110 10124
rect 18104 10115 18132 10121
rect 18120 10081 18132 10115
rect 18104 10075 18132 10081
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10112 18291 10115
rect 18966 10112 18972 10124
rect 18279 10084 18972 10112
rect 18279 10081 18291 10084
rect 18233 10075 18291 10081
rect 18104 10072 18110 10075
rect 18966 10072 18972 10084
rect 19024 10072 19030 10124
rect 21266 10112 21272 10124
rect 21227 10084 21272 10112
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21542 10112 21548 10124
rect 21503 10084 21548 10112
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10013 17095 10047
rect 19426 10044 19432 10056
rect 19387 10016 19432 10044
rect 17037 10007 17095 10013
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 16577 9911 16635 9917
rect 16577 9908 16589 9911
rect 2556 9880 16589 9908
rect 2556 9868 2562 9880
rect 16577 9877 16589 9880
rect 16623 9908 16635 9911
rect 16850 9908 16856 9920
rect 16623 9880 16856 9908
rect 16623 9877 16635 9880
rect 16577 9871 16635 9877
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 17052 9908 17080 10007
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 19702 10044 19708 10056
rect 19663 10016 19708 10044
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 19978 9976 19984 9988
rect 18708 9948 19984 9976
rect 17678 9908 17684 9920
rect 17052 9880 17684 9908
rect 17678 9868 17684 9880
rect 17736 9908 17742 9920
rect 18708 9908 18736 9948
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 18874 9908 18880 9920
rect 17736 9880 18736 9908
rect 18835 9880 18880 9908
rect 17736 9868 17742 9880
rect 18874 9868 18880 9880
rect 18932 9868 18938 9920
rect 1104 9818 22976 9840
rect 1104 9766 6378 9818
rect 6430 9766 6442 9818
rect 6494 9766 6506 9818
rect 6558 9766 6570 9818
rect 6622 9766 6634 9818
rect 6686 9766 11806 9818
rect 11858 9766 11870 9818
rect 11922 9766 11934 9818
rect 11986 9766 11998 9818
rect 12050 9766 12062 9818
rect 12114 9766 17234 9818
rect 17286 9766 17298 9818
rect 17350 9766 17362 9818
rect 17414 9766 17426 9818
rect 17478 9766 17490 9818
rect 17542 9766 22662 9818
rect 22714 9766 22726 9818
rect 22778 9766 22790 9818
rect 22842 9766 22854 9818
rect 22906 9766 22918 9818
rect 22970 9766 22976 9818
rect 1104 9744 22976 9766
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18141 9707 18199 9713
rect 18141 9704 18153 9707
rect 18104 9676 18153 9704
rect 18104 9664 18110 9676
rect 18141 9673 18153 9676
rect 18187 9673 18199 9707
rect 18141 9667 18199 9673
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 18785 9707 18843 9713
rect 18785 9704 18797 9707
rect 18656 9676 18797 9704
rect 18656 9664 18662 9676
rect 18785 9673 18797 9676
rect 18831 9673 18843 9707
rect 19426 9704 19432 9716
rect 19387 9676 19432 9704
rect 18785 9667 18843 9673
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 19978 9704 19984 9716
rect 19939 9676 19984 9704
rect 19978 9664 19984 9676
rect 20036 9664 20042 9716
rect 21358 9636 21364 9648
rect 21008 9608 21364 9636
rect 18690 9568 18696 9580
rect 18651 9540 18696 9568
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 18892 9500 18920 9531
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 21008 9577 21036 9608
rect 21358 9596 21364 9608
rect 21416 9596 21422 9648
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 19300 9540 19349 9568
rect 19300 9528 19306 9540
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 19337 9531 19395 9537
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9537 21051 9571
rect 21174 9568 21180 9580
rect 21135 9540 21180 9568
rect 20993 9531 21051 9537
rect 19536 9500 19564 9531
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 20346 9500 20352 9512
rect 18892 9472 20352 9500
rect 20346 9460 20352 9472
rect 20404 9500 20410 9512
rect 21085 9503 21143 9509
rect 21085 9500 21097 9503
rect 20404 9472 21097 9500
rect 20404 9460 20410 9472
rect 21085 9469 21097 9472
rect 21131 9469 21143 9503
rect 21085 9463 21143 9469
rect 1104 9274 22816 9296
rect 1104 9222 3664 9274
rect 3716 9222 3728 9274
rect 3780 9222 3792 9274
rect 3844 9222 3856 9274
rect 3908 9222 3920 9274
rect 3972 9222 9092 9274
rect 9144 9222 9156 9274
rect 9208 9222 9220 9274
rect 9272 9222 9284 9274
rect 9336 9222 9348 9274
rect 9400 9222 14520 9274
rect 14572 9222 14584 9274
rect 14636 9222 14648 9274
rect 14700 9222 14712 9274
rect 14764 9222 14776 9274
rect 14828 9222 19948 9274
rect 20000 9222 20012 9274
rect 20064 9222 20076 9274
rect 20128 9222 20140 9274
rect 20192 9222 20204 9274
rect 20256 9222 22816 9274
rect 1104 9200 22816 9222
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 21634 8820 21640 8832
rect 20588 8792 21640 8820
rect 20588 8780 20594 8792
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 1104 8730 22976 8752
rect 1104 8678 6378 8730
rect 6430 8678 6442 8730
rect 6494 8678 6506 8730
rect 6558 8678 6570 8730
rect 6622 8678 6634 8730
rect 6686 8678 11806 8730
rect 11858 8678 11870 8730
rect 11922 8678 11934 8730
rect 11986 8678 11998 8730
rect 12050 8678 12062 8730
rect 12114 8678 17234 8730
rect 17286 8678 17298 8730
rect 17350 8678 17362 8730
rect 17414 8678 17426 8730
rect 17478 8678 17490 8730
rect 17542 8678 22662 8730
rect 22714 8678 22726 8730
rect 22778 8678 22790 8730
rect 22842 8678 22854 8730
rect 22906 8678 22918 8730
rect 22970 8678 22976 8730
rect 1104 8656 22976 8678
rect 19168 8588 19334 8616
rect 19168 8492 19196 8588
rect 19306 8548 19334 8588
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 21692 8588 22048 8616
rect 21692 8576 21698 8588
rect 22020 8557 22048 8588
rect 22005 8551 22063 8557
rect 19306 8520 21312 8548
rect 19150 8480 19156 8492
rect 19111 8452 19156 8480
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 20346 8480 20352 8492
rect 20303 8452 20352 8480
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 20530 8372 20536 8424
rect 20588 8412 20594 8424
rect 20588 8384 20633 8412
rect 20588 8372 20594 8384
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 18693 8347 18751 8353
rect 18693 8344 18705 8347
rect 18656 8316 18705 8344
rect 18656 8304 18662 8316
rect 18693 8313 18705 8316
rect 18739 8313 18751 8347
rect 18693 8307 18751 8313
rect 20349 8347 20407 8353
rect 20349 8313 20361 8347
rect 20395 8344 20407 8347
rect 20990 8344 20996 8356
rect 20395 8316 20852 8344
rect 20951 8316 20996 8344
rect 20395 8313 20407 8316
rect 20349 8307 20407 8313
rect 18874 8276 18880 8288
rect 18835 8248 18880 8276
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 20438 8276 20444 8288
rect 20399 8248 20444 8276
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 20824 8276 20852 8316
rect 20990 8304 20996 8316
rect 21048 8304 21054 8356
rect 21192 8344 21220 8443
rect 21284 8412 21312 8520
rect 22005 8517 22017 8551
rect 22051 8517 22063 8551
rect 22005 8511 22063 8517
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 21284 8384 21465 8412
rect 21453 8381 21465 8384
rect 21499 8412 21511 8415
rect 22204 8412 22232 8443
rect 21499 8384 22232 8412
rect 21499 8381 21511 8384
rect 21453 8375 21511 8381
rect 22005 8347 22063 8353
rect 22005 8344 22017 8347
rect 21192 8316 22017 8344
rect 22005 8313 22017 8316
rect 22051 8313 22063 8347
rect 22005 8307 22063 8313
rect 21361 8279 21419 8285
rect 21361 8276 21373 8279
rect 20824 8248 21373 8276
rect 21361 8245 21373 8248
rect 21407 8276 21419 8279
rect 21542 8276 21548 8288
rect 21407 8248 21548 8276
rect 21407 8245 21419 8248
rect 21361 8239 21419 8245
rect 21542 8236 21548 8248
rect 21600 8276 21606 8288
rect 22296 8276 22324 8443
rect 21600 8248 22324 8276
rect 21600 8236 21606 8248
rect 1104 8186 22816 8208
rect 1104 8134 3664 8186
rect 3716 8134 3728 8186
rect 3780 8134 3792 8186
rect 3844 8134 3856 8186
rect 3908 8134 3920 8186
rect 3972 8134 9092 8186
rect 9144 8134 9156 8186
rect 9208 8134 9220 8186
rect 9272 8134 9284 8186
rect 9336 8134 9348 8186
rect 9400 8134 14520 8186
rect 14572 8134 14584 8186
rect 14636 8134 14648 8186
rect 14700 8134 14712 8186
rect 14764 8134 14776 8186
rect 14828 8134 19948 8186
rect 20000 8134 20012 8186
rect 20064 8134 20076 8186
rect 20128 8134 20140 8186
rect 20192 8134 20204 8186
rect 20256 8134 22816 8186
rect 1104 8112 22816 8134
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 18196 7908 19472 7936
rect 18196 7896 18202 7908
rect 18046 7868 18052 7880
rect 18007 7840 18052 7868
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18414 7868 18420 7880
rect 18375 7840 18420 7868
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18874 7868 18880 7880
rect 18835 7840 18880 7868
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19444 7877 19472 7908
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 18601 7803 18659 7809
rect 18601 7769 18613 7803
rect 18647 7800 18659 7803
rect 18690 7800 18696 7812
rect 18647 7772 18696 7800
rect 18647 7769 18659 7772
rect 18601 7763 18659 7769
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 18892 7800 18920 7828
rect 19150 7800 19156 7812
rect 18892 7772 19156 7800
rect 19150 7760 19156 7772
rect 19208 7800 19214 7812
rect 19613 7803 19671 7809
rect 19613 7800 19625 7803
rect 19208 7772 19625 7800
rect 19208 7760 19214 7772
rect 19613 7769 19625 7772
rect 19659 7769 19671 7803
rect 19613 7763 19671 7769
rect 18506 7692 18512 7744
rect 18564 7732 18570 7744
rect 19797 7735 19855 7741
rect 19797 7732 19809 7735
rect 18564 7704 19809 7732
rect 18564 7692 18570 7704
rect 19797 7701 19809 7704
rect 19843 7701 19855 7735
rect 19797 7695 19855 7701
rect 1104 7642 22976 7664
rect 1104 7590 6378 7642
rect 6430 7590 6442 7642
rect 6494 7590 6506 7642
rect 6558 7590 6570 7642
rect 6622 7590 6634 7642
rect 6686 7590 11806 7642
rect 11858 7590 11870 7642
rect 11922 7590 11934 7642
rect 11986 7590 11998 7642
rect 12050 7590 12062 7642
rect 12114 7590 17234 7642
rect 17286 7590 17298 7642
rect 17350 7590 17362 7642
rect 17414 7590 17426 7642
rect 17478 7590 17490 7642
rect 17542 7590 22662 7642
rect 22714 7590 22726 7642
rect 22778 7590 22790 7642
rect 22842 7590 22854 7642
rect 22906 7590 22918 7642
rect 22970 7590 22976 7642
rect 1104 7568 22976 7590
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7528 18843 7531
rect 19242 7528 19248 7540
rect 18831 7500 19248 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 20530 7460 20536 7472
rect 18104 7432 20536 7460
rect 18104 7420 18110 7432
rect 18616 7401 18644 7432
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 18601 7395 18659 7401
rect 18601 7361 18613 7395
rect 18647 7361 18659 7395
rect 18874 7392 18880 7404
rect 18835 7364 18880 7392
rect 18601 7355 18659 7361
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 18414 7324 18420 7336
rect 18375 7296 18420 7324
rect 18414 7284 18420 7296
rect 18472 7284 18478 7336
rect 1104 7098 22816 7120
rect 1104 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 9092 7098
rect 9144 7046 9156 7098
rect 9208 7046 9220 7098
rect 9272 7046 9284 7098
rect 9336 7046 9348 7098
rect 9400 7046 14520 7098
rect 14572 7046 14584 7098
rect 14636 7046 14648 7098
rect 14700 7046 14712 7098
rect 14764 7046 14776 7098
rect 14828 7046 19948 7098
rect 20000 7046 20012 7098
rect 20064 7046 20076 7098
rect 20128 7046 20140 7098
rect 20192 7046 20204 7098
rect 20256 7046 22816 7098
rect 1104 7024 22816 7046
rect 1104 6554 22976 6576
rect 1104 6502 6378 6554
rect 6430 6502 6442 6554
rect 6494 6502 6506 6554
rect 6558 6502 6570 6554
rect 6622 6502 6634 6554
rect 6686 6502 11806 6554
rect 11858 6502 11870 6554
rect 11922 6502 11934 6554
rect 11986 6502 11998 6554
rect 12050 6502 12062 6554
rect 12114 6502 17234 6554
rect 17286 6502 17298 6554
rect 17350 6502 17362 6554
rect 17414 6502 17426 6554
rect 17478 6502 17490 6554
rect 17542 6502 22662 6554
rect 22714 6502 22726 6554
rect 22778 6502 22790 6554
rect 22842 6502 22854 6554
rect 22906 6502 22918 6554
rect 22970 6502 22976 6554
rect 1104 6480 22976 6502
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 21453 6443 21511 6449
rect 21453 6440 21465 6443
rect 21232 6412 21465 6440
rect 21232 6400 21238 6412
rect 21453 6409 21465 6412
rect 21499 6409 21511 6443
rect 21453 6403 21511 6409
rect 20340 6375 20398 6381
rect 20340 6341 20352 6375
rect 20386 6372 20398 6375
rect 20438 6372 20444 6384
rect 20386 6344 20444 6372
rect 20386 6341 20398 6344
rect 20340 6335 20398 6341
rect 20438 6332 20444 6344
rect 20496 6332 20502 6384
rect 20073 6239 20131 6245
rect 20073 6205 20085 6239
rect 20119 6205 20131 6239
rect 20073 6199 20131 6205
rect 20088 6100 20116 6199
rect 20438 6100 20444 6112
rect 20088 6072 20444 6100
rect 20438 6060 20444 6072
rect 20496 6060 20502 6112
rect 1104 6010 22816 6032
rect 1104 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 9092 6010
rect 9144 5958 9156 6010
rect 9208 5958 9220 6010
rect 9272 5958 9284 6010
rect 9336 5958 9348 6010
rect 9400 5958 14520 6010
rect 14572 5958 14584 6010
rect 14636 5958 14648 6010
rect 14700 5958 14712 6010
rect 14764 5958 14776 6010
rect 14828 5958 19948 6010
rect 20000 5958 20012 6010
rect 20064 5958 20076 6010
rect 20128 5958 20140 6010
rect 20192 5958 20204 6010
rect 20256 5958 22816 6010
rect 1104 5936 22816 5958
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 20073 5695 20131 5701
rect 20073 5692 20085 5695
rect 19392 5664 20085 5692
rect 19392 5652 19398 5664
rect 20073 5661 20085 5664
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 19610 5584 19616 5636
rect 19668 5624 19674 5636
rect 20318 5627 20376 5633
rect 20318 5624 20330 5627
rect 19668 5596 20330 5624
rect 19668 5584 19674 5596
rect 20318 5593 20330 5596
rect 20364 5593 20376 5627
rect 20318 5587 20376 5593
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 21453 5559 21511 5565
rect 21453 5556 21465 5559
rect 18288 5528 21465 5556
rect 18288 5516 18294 5528
rect 21453 5525 21465 5528
rect 21499 5525 21511 5559
rect 21453 5519 21511 5525
rect 1104 5466 22976 5488
rect 1104 5414 6378 5466
rect 6430 5414 6442 5466
rect 6494 5414 6506 5466
rect 6558 5414 6570 5466
rect 6622 5414 6634 5466
rect 6686 5414 11806 5466
rect 11858 5414 11870 5466
rect 11922 5414 11934 5466
rect 11986 5414 11998 5466
rect 12050 5414 12062 5466
rect 12114 5414 17234 5466
rect 17286 5414 17298 5466
rect 17350 5414 17362 5466
rect 17414 5414 17426 5466
rect 17478 5414 17490 5466
rect 17542 5414 22662 5466
rect 22714 5414 22726 5466
rect 22778 5414 22790 5466
rect 22842 5414 22854 5466
rect 22906 5414 22918 5466
rect 22970 5414 22976 5466
rect 1104 5392 22976 5414
rect 20438 5312 20444 5364
rect 20496 5352 20502 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 20496 5324 20637 5352
rect 20496 5312 20502 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 19981 5287 20039 5293
rect 19981 5253 19993 5287
rect 20027 5284 20039 5287
rect 20806 5284 20812 5296
rect 20027 5256 20812 5284
rect 20027 5253 20039 5256
rect 19981 5247 20039 5253
rect 20806 5244 20812 5256
rect 20864 5244 20870 5296
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 19392 5188 20545 5216
rect 19392 5176 19398 5188
rect 20533 5185 20545 5188
rect 20579 5185 20591 5219
rect 20533 5179 20591 5185
rect 18693 5015 18751 5021
rect 18693 4981 18705 5015
rect 18739 5012 18751 5015
rect 19334 5012 19340 5024
rect 18739 4984 19340 5012
rect 18739 4981 18751 4984
rect 18693 4975 18751 4981
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 1104 4922 22816 4944
rect 1104 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 9092 4922
rect 9144 4870 9156 4922
rect 9208 4870 9220 4922
rect 9272 4870 9284 4922
rect 9336 4870 9348 4922
rect 9400 4870 14520 4922
rect 14572 4870 14584 4922
rect 14636 4870 14648 4922
rect 14700 4870 14712 4922
rect 14764 4870 14776 4922
rect 14828 4870 19948 4922
rect 20000 4870 20012 4922
rect 20064 4870 20076 4922
rect 20128 4870 20140 4922
rect 20192 4870 20204 4922
rect 20256 4870 22816 4922
rect 1104 4848 22816 4870
rect 18877 4811 18935 4817
rect 18877 4777 18889 4811
rect 18923 4808 18935 4811
rect 19610 4808 19616 4820
rect 18923 4780 19616 4808
rect 18923 4777 18935 4780
rect 18877 4771 18935 4777
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 20257 4811 20315 4817
rect 20257 4777 20269 4811
rect 20303 4808 20315 4811
rect 20530 4808 20536 4820
rect 20303 4780 20536 4808
rect 20303 4777 20315 4780
rect 20257 4771 20315 4777
rect 15654 4700 15660 4752
rect 15712 4740 15718 4752
rect 15712 4712 19334 4740
rect 15712 4700 15718 4712
rect 18230 4672 18236 4684
rect 18191 4644 18236 4672
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 18432 4613 18460 4712
rect 19306 4672 19334 4712
rect 19306 4644 19472 4672
rect 18391 4607 18460 4613
rect 18391 4573 18403 4607
rect 18437 4576 18460 4607
rect 18598 4604 18604 4616
rect 18559 4576 18604 4604
rect 18437 4573 18449 4576
rect 18391 4567 18449 4573
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 19444 4613 19472 4644
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4573 18751 4607
rect 18693 4567 18751 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 18506 4496 18512 4548
rect 18564 4536 18570 4548
rect 18708 4536 18736 4567
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 20272 4604 20300 4771
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 19668 4576 20300 4604
rect 21637 4607 21695 4613
rect 19668 4564 19674 4576
rect 21637 4573 21649 4607
rect 21683 4604 21695 4607
rect 22094 4604 22100 4616
rect 21683 4576 22100 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 22094 4564 22100 4576
rect 22152 4564 22158 4616
rect 19521 4539 19579 4545
rect 19521 4536 19533 4539
rect 18564 4508 18609 4536
rect 18708 4508 19533 4536
rect 18564 4496 18570 4508
rect 19521 4505 19533 4508
rect 19567 4505 19579 4539
rect 19521 4499 19579 4505
rect 21392 4539 21450 4545
rect 21392 4505 21404 4539
rect 21438 4536 21450 4539
rect 22002 4536 22008 4548
rect 21438 4508 22008 4536
rect 21438 4505 21450 4508
rect 21392 4499 21450 4505
rect 22002 4496 22008 4508
rect 22060 4496 22066 4548
rect 22186 4468 22192 4480
rect 22147 4440 22192 4468
rect 22186 4428 22192 4440
rect 22244 4428 22250 4480
rect 1104 4378 22976 4400
rect 1104 4326 6378 4378
rect 6430 4326 6442 4378
rect 6494 4326 6506 4378
rect 6558 4326 6570 4378
rect 6622 4326 6634 4378
rect 6686 4326 11806 4378
rect 11858 4326 11870 4378
rect 11922 4326 11934 4378
rect 11986 4326 11998 4378
rect 12050 4326 12062 4378
rect 12114 4326 17234 4378
rect 17286 4326 17298 4378
rect 17350 4326 17362 4378
rect 17414 4326 17426 4378
rect 17478 4326 17490 4378
rect 17542 4326 22662 4378
rect 22714 4326 22726 4378
rect 22778 4326 22790 4378
rect 22842 4326 22854 4378
rect 22906 4326 22918 4378
rect 22970 4326 22976 4378
rect 1104 4304 22976 4326
rect 19334 4128 19340 4140
rect 19295 4100 19340 4128
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 20237 4131 20295 4137
rect 20237 4128 20249 4131
rect 19576 4100 20249 4128
rect 19576 4088 19582 4100
rect 20237 4097 20249 4100
rect 20283 4097 20295 4131
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 20237 4091 20295 4097
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 19429 4063 19487 4069
rect 19429 4029 19441 4063
rect 19475 4060 19487 4063
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19475 4032 19993 4060
rect 19475 4029 19487 4032
rect 19429 4023 19487 4029
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 21358 3924 21364 3936
rect 21319 3896 21364 3924
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 1104 3834 22816 3856
rect 1104 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 9092 3834
rect 9144 3782 9156 3834
rect 9208 3782 9220 3834
rect 9272 3782 9284 3834
rect 9336 3782 9348 3834
rect 9400 3782 14520 3834
rect 14572 3782 14584 3834
rect 14636 3782 14648 3834
rect 14700 3782 14712 3834
rect 14764 3782 14776 3834
rect 14828 3782 19948 3834
rect 20000 3782 20012 3834
rect 20064 3782 20076 3834
rect 20128 3782 20140 3834
rect 20192 3782 20204 3834
rect 20256 3782 22816 3834
rect 1104 3760 22816 3782
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 19518 3720 19524 3732
rect 18371 3692 19524 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 20806 3720 20812 3732
rect 20767 3692 20812 3720
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21358 3584 21364 3596
rect 18156 3556 21364 3584
rect 18156 3525 18184 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 19610 3516 19616 3528
rect 18371 3488 19616 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 22186 3448 22192 3460
rect 21876 3420 22192 3448
rect 21876 3408 21882 3420
rect 22186 3408 22192 3420
rect 22244 3448 22250 3460
rect 22281 3451 22339 3457
rect 22281 3448 22293 3451
rect 22244 3420 22293 3448
rect 22244 3408 22250 3420
rect 22281 3417 22293 3420
rect 22327 3417 22339 3451
rect 22281 3411 22339 3417
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 14366 3380 14372 3392
rect 13044 3352 14372 3380
rect 13044 3340 13050 3352
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 1104 3290 22976 3312
rect 1104 3238 6378 3290
rect 6430 3238 6442 3290
rect 6494 3238 6506 3290
rect 6558 3238 6570 3290
rect 6622 3238 6634 3290
rect 6686 3238 11806 3290
rect 11858 3238 11870 3290
rect 11922 3238 11934 3290
rect 11986 3238 11998 3290
rect 12050 3238 12062 3290
rect 12114 3238 17234 3290
rect 17286 3238 17298 3290
rect 17350 3238 17362 3290
rect 17414 3238 17426 3290
rect 17478 3238 17490 3290
rect 17542 3238 22662 3290
rect 22714 3238 22726 3290
rect 22778 3238 22790 3290
rect 22842 3238 22854 3290
rect 22906 3238 22918 3290
rect 22970 3238 22976 3290
rect 1104 3216 22976 3238
rect 13173 3179 13231 3185
rect 13173 3145 13185 3179
rect 13219 3176 13231 3179
rect 18414 3176 18420 3188
rect 13219 3148 18420 3176
rect 13219 3145 13231 3148
rect 13173 3139 13231 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 22094 3176 22100 3188
rect 22055 3148 22100 3176
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 18230 3108 18236 3120
rect 13372 3080 14320 3108
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13372 3049 13400 3080
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 14090 3040 14096 3052
rect 13679 3012 14096 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 13372 2972 13400 3003
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 12400 2944 13400 2972
rect 14185 2975 14243 2981
rect 12400 2932 12406 2944
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14200 2904 14228 2935
rect 13464 2876 14228 2904
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 13464 2845 13492 2876
rect 14292 2845 14320 3080
rect 17880 3080 18236 3108
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 17880 3049 17908 3080
rect 18230 3068 18236 3080
rect 18288 3068 18294 3120
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 14424 3012 15577 3040
rect 14424 3000 14430 3012
rect 15565 3009 15577 3012
rect 15611 3009 15623 3043
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 15565 3003 15623 3009
rect 15764 3012 16865 3040
rect 14553 2907 14611 2913
rect 14553 2873 14565 2907
rect 14599 2904 14611 2907
rect 15654 2904 15660 2916
rect 14599 2876 15660 2904
rect 14599 2873 14611 2876
rect 14553 2867 14611 2873
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 15764 2913 15792 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3009 17923 3043
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 17865 3003 17923 3009
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 19702 2972 19708 2984
rect 18371 2944 19708 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 15749 2907 15807 2913
rect 15749 2873 15761 2907
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 17037 2907 17095 2913
rect 17037 2873 17049 2907
rect 17083 2904 17095 2907
rect 18064 2904 18092 2935
rect 17083 2876 18092 2904
rect 17083 2873 17095 2876
rect 17037 2867 17095 2873
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 13412 2808 13461 2836
rect 13412 2796 13418 2808
rect 13449 2805 13461 2808
rect 13495 2805 13507 2839
rect 13449 2799 13507 2805
rect 14277 2839 14335 2845
rect 14277 2805 14289 2839
rect 14323 2805 14335 2839
rect 14277 2799 14335 2805
rect 17862 2796 17868 2848
rect 17920 2836 17926 2848
rect 18340 2836 18368 2935
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 17920 2808 18368 2836
rect 17920 2796 17926 2808
rect 1104 2746 22816 2768
rect 1104 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 9092 2746
rect 9144 2694 9156 2746
rect 9208 2694 9220 2746
rect 9272 2694 9284 2746
rect 9336 2694 9348 2746
rect 9400 2694 14520 2746
rect 14572 2694 14584 2746
rect 14636 2694 14648 2746
rect 14700 2694 14712 2746
rect 14764 2694 14776 2746
rect 14828 2694 19948 2746
rect 20000 2694 20012 2746
rect 20064 2694 20076 2746
rect 20128 2694 20140 2746
rect 20192 2694 20204 2746
rect 20256 2694 22816 2746
rect 1104 2672 22816 2694
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 12342 2632 12348 2644
rect 10275 2604 12348 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14090 2592 14096 2644
rect 14148 2632 14154 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 14148 2604 14289 2632
rect 14148 2592 14154 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 17497 2635 17555 2641
rect 17497 2601 17509 2635
rect 17543 2632 17555 2635
rect 18874 2632 18880 2644
rect 17543 2604 18880 2632
rect 17543 2601 17555 2604
rect 17497 2595 17555 2601
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 12986 2564 12992 2576
rect 2363 2536 12992 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 22097 2499 22155 2505
rect 22097 2496 22109 2499
rect 18923 2468 22109 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 22097 2465 22109 2468
rect 22143 2465 22155 2499
rect 22097 2459 22155 2465
rect 2038 2388 2044 2440
rect 2096 2428 2102 2440
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 2096 2400 2145 2428
rect 2096 2388 2102 2400
rect 2133 2397 2145 2400
rect 2179 2428 2191 2431
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2179 2400 2789 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6052 2400 6561 2428
rect 6052 2388 6058 2400
rect 6549 2397 6561 2400
rect 6595 2428 6607 2431
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6595 2400 7205 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 10008 2400 10057 2428
rect 10008 2388 10014 2400
rect 10045 2397 10057 2400
rect 10091 2428 10103 2431
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10091 2400 10701 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13964 2400 14473 2428
rect 13964 2388 13970 2400
rect 14461 2397 14473 2400
rect 14507 2428 14519 2431
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14507 2400 14933 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 19705 2431 19763 2437
rect 19705 2397 19717 2431
rect 19751 2428 19763 2431
rect 20806 2428 20812 2440
rect 19751 2400 20812 2428
rect 19751 2397 19763 2400
rect 19705 2391 19763 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2428 21511 2431
rect 22002 2428 22008 2440
rect 21499 2400 22008 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 18632 2363 18690 2369
rect 18632 2329 18644 2363
rect 18678 2360 18690 2363
rect 20990 2360 20996 2372
rect 18678 2332 20996 2360
rect 18678 2329 18690 2332
rect 18632 2323 18690 2329
rect 20990 2320 20996 2332
rect 21048 2320 21054 2372
rect 6733 2295 6791 2301
rect 6733 2261 6745 2295
rect 6779 2292 6791 2295
rect 13354 2292 13360 2304
rect 6779 2264 13360 2292
rect 6779 2261 6791 2264
rect 6733 2255 6791 2261
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 1104 2202 22976 2224
rect 1104 2150 6378 2202
rect 6430 2150 6442 2202
rect 6494 2150 6506 2202
rect 6558 2150 6570 2202
rect 6622 2150 6634 2202
rect 6686 2150 11806 2202
rect 11858 2150 11870 2202
rect 11922 2150 11934 2202
rect 11986 2150 11998 2202
rect 12050 2150 12062 2202
rect 12114 2150 17234 2202
rect 17286 2150 17298 2202
rect 17350 2150 17362 2202
rect 17414 2150 17426 2202
rect 17478 2150 17490 2202
rect 17542 2150 22662 2202
rect 22714 2150 22726 2202
rect 22778 2150 22790 2202
rect 22842 2150 22854 2202
rect 22906 2150 22918 2202
rect 22970 2150 22976 2202
rect 1104 2128 22976 2150
<< via1 >>
rect 6378 21734 6430 21786
rect 6442 21734 6494 21786
rect 6506 21734 6558 21786
rect 6570 21734 6622 21786
rect 6634 21734 6686 21786
rect 11806 21734 11858 21786
rect 11870 21734 11922 21786
rect 11934 21734 11986 21786
rect 11998 21734 12050 21786
rect 12062 21734 12114 21786
rect 17234 21734 17286 21786
rect 17298 21734 17350 21786
rect 17362 21734 17414 21786
rect 17426 21734 17478 21786
rect 17490 21734 17542 21786
rect 22662 21734 22714 21786
rect 22726 21734 22778 21786
rect 22790 21734 22842 21786
rect 22854 21734 22906 21786
rect 22918 21734 22970 21786
rect 1860 21675 1912 21684
rect 1860 21641 1869 21675
rect 1869 21641 1903 21675
rect 1903 21641 1912 21675
rect 1860 21632 1912 21641
rect 4804 21675 4856 21684
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 7748 21675 7800 21684
rect 7748 21641 7757 21675
rect 7757 21641 7791 21675
rect 7791 21641 7800 21675
rect 7748 21632 7800 21641
rect 10692 21675 10744 21684
rect 10692 21641 10701 21675
rect 10701 21641 10735 21675
rect 10735 21641 10744 21675
rect 10692 21632 10744 21641
rect 13820 21632 13872 21684
rect 16580 21632 16632 21684
rect 19524 21675 19576 21684
rect 19524 21641 19533 21675
rect 19533 21641 19567 21675
rect 19567 21641 19576 21675
rect 19524 21632 19576 21641
rect 22192 21675 22244 21684
rect 22192 21641 22201 21675
rect 22201 21641 22235 21675
rect 22235 21641 22244 21675
rect 22192 21632 22244 21641
rect 2504 21496 2556 21548
rect 2504 21335 2556 21344
rect 2504 21301 2513 21335
rect 2513 21301 2547 21335
rect 2547 21301 2556 21335
rect 2504 21292 2556 21301
rect 8392 21496 8444 21548
rect 11704 21496 11756 21548
rect 17868 21496 17920 21548
rect 20444 21496 20496 21548
rect 19064 21428 19116 21480
rect 19800 21428 19852 21480
rect 6184 21292 6236 21344
rect 8392 21335 8444 21344
rect 8392 21301 8401 21335
rect 8401 21301 8435 21335
rect 8435 21301 8444 21335
rect 8392 21292 8444 21301
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 3664 21190 3716 21242
rect 3728 21190 3780 21242
rect 3792 21190 3844 21242
rect 3856 21190 3908 21242
rect 3920 21190 3972 21242
rect 9092 21190 9144 21242
rect 9156 21190 9208 21242
rect 9220 21190 9272 21242
rect 9284 21190 9336 21242
rect 9348 21190 9400 21242
rect 14520 21190 14572 21242
rect 14584 21190 14636 21242
rect 14648 21190 14700 21242
rect 14712 21190 14764 21242
rect 14776 21190 14828 21242
rect 19948 21190 20000 21242
rect 20012 21190 20064 21242
rect 20076 21190 20128 21242
rect 20140 21190 20192 21242
rect 20204 21190 20256 21242
rect 6378 20646 6430 20698
rect 6442 20646 6494 20698
rect 6506 20646 6558 20698
rect 6570 20646 6622 20698
rect 6634 20646 6686 20698
rect 11806 20646 11858 20698
rect 11870 20646 11922 20698
rect 11934 20646 11986 20698
rect 11998 20646 12050 20698
rect 12062 20646 12114 20698
rect 17234 20646 17286 20698
rect 17298 20646 17350 20698
rect 17362 20646 17414 20698
rect 17426 20646 17478 20698
rect 17490 20646 17542 20698
rect 22662 20646 22714 20698
rect 22726 20646 22778 20698
rect 22790 20646 22842 20698
rect 22854 20646 22906 20698
rect 22918 20646 22970 20698
rect 3664 20102 3716 20154
rect 3728 20102 3780 20154
rect 3792 20102 3844 20154
rect 3856 20102 3908 20154
rect 3920 20102 3972 20154
rect 9092 20102 9144 20154
rect 9156 20102 9208 20154
rect 9220 20102 9272 20154
rect 9284 20102 9336 20154
rect 9348 20102 9400 20154
rect 14520 20102 14572 20154
rect 14584 20102 14636 20154
rect 14648 20102 14700 20154
rect 14712 20102 14764 20154
rect 14776 20102 14828 20154
rect 19948 20102 20000 20154
rect 20012 20102 20064 20154
rect 20076 20102 20128 20154
rect 20140 20102 20192 20154
rect 20204 20102 20256 20154
rect 6378 19558 6430 19610
rect 6442 19558 6494 19610
rect 6506 19558 6558 19610
rect 6570 19558 6622 19610
rect 6634 19558 6686 19610
rect 11806 19558 11858 19610
rect 11870 19558 11922 19610
rect 11934 19558 11986 19610
rect 11998 19558 12050 19610
rect 12062 19558 12114 19610
rect 17234 19558 17286 19610
rect 17298 19558 17350 19610
rect 17362 19558 17414 19610
rect 17426 19558 17478 19610
rect 17490 19558 17542 19610
rect 22662 19558 22714 19610
rect 22726 19558 22778 19610
rect 22790 19558 22842 19610
rect 22854 19558 22906 19610
rect 22918 19558 22970 19610
rect 3664 19014 3716 19066
rect 3728 19014 3780 19066
rect 3792 19014 3844 19066
rect 3856 19014 3908 19066
rect 3920 19014 3972 19066
rect 9092 19014 9144 19066
rect 9156 19014 9208 19066
rect 9220 19014 9272 19066
rect 9284 19014 9336 19066
rect 9348 19014 9400 19066
rect 14520 19014 14572 19066
rect 14584 19014 14636 19066
rect 14648 19014 14700 19066
rect 14712 19014 14764 19066
rect 14776 19014 14828 19066
rect 19948 19014 20000 19066
rect 20012 19014 20064 19066
rect 20076 19014 20128 19066
rect 20140 19014 20192 19066
rect 20204 19014 20256 19066
rect 6378 18470 6430 18522
rect 6442 18470 6494 18522
rect 6506 18470 6558 18522
rect 6570 18470 6622 18522
rect 6634 18470 6686 18522
rect 11806 18470 11858 18522
rect 11870 18470 11922 18522
rect 11934 18470 11986 18522
rect 11998 18470 12050 18522
rect 12062 18470 12114 18522
rect 17234 18470 17286 18522
rect 17298 18470 17350 18522
rect 17362 18470 17414 18522
rect 17426 18470 17478 18522
rect 17490 18470 17542 18522
rect 22662 18470 22714 18522
rect 22726 18470 22778 18522
rect 22790 18470 22842 18522
rect 22854 18470 22906 18522
rect 22918 18470 22970 18522
rect 3664 17926 3716 17978
rect 3728 17926 3780 17978
rect 3792 17926 3844 17978
rect 3856 17926 3908 17978
rect 3920 17926 3972 17978
rect 9092 17926 9144 17978
rect 9156 17926 9208 17978
rect 9220 17926 9272 17978
rect 9284 17926 9336 17978
rect 9348 17926 9400 17978
rect 14520 17926 14572 17978
rect 14584 17926 14636 17978
rect 14648 17926 14700 17978
rect 14712 17926 14764 17978
rect 14776 17926 14828 17978
rect 19948 17926 20000 17978
rect 20012 17926 20064 17978
rect 20076 17926 20128 17978
rect 20140 17926 20192 17978
rect 20204 17926 20256 17978
rect 6378 17382 6430 17434
rect 6442 17382 6494 17434
rect 6506 17382 6558 17434
rect 6570 17382 6622 17434
rect 6634 17382 6686 17434
rect 11806 17382 11858 17434
rect 11870 17382 11922 17434
rect 11934 17382 11986 17434
rect 11998 17382 12050 17434
rect 12062 17382 12114 17434
rect 17234 17382 17286 17434
rect 17298 17382 17350 17434
rect 17362 17382 17414 17434
rect 17426 17382 17478 17434
rect 17490 17382 17542 17434
rect 22662 17382 22714 17434
rect 22726 17382 22778 17434
rect 22790 17382 22842 17434
rect 22854 17382 22906 17434
rect 22918 17382 22970 17434
rect 3664 16838 3716 16890
rect 3728 16838 3780 16890
rect 3792 16838 3844 16890
rect 3856 16838 3908 16890
rect 3920 16838 3972 16890
rect 9092 16838 9144 16890
rect 9156 16838 9208 16890
rect 9220 16838 9272 16890
rect 9284 16838 9336 16890
rect 9348 16838 9400 16890
rect 14520 16838 14572 16890
rect 14584 16838 14636 16890
rect 14648 16838 14700 16890
rect 14712 16838 14764 16890
rect 14776 16838 14828 16890
rect 19948 16838 20000 16890
rect 20012 16838 20064 16890
rect 20076 16838 20128 16890
rect 20140 16838 20192 16890
rect 20204 16838 20256 16890
rect 6378 16294 6430 16346
rect 6442 16294 6494 16346
rect 6506 16294 6558 16346
rect 6570 16294 6622 16346
rect 6634 16294 6686 16346
rect 11806 16294 11858 16346
rect 11870 16294 11922 16346
rect 11934 16294 11986 16346
rect 11998 16294 12050 16346
rect 12062 16294 12114 16346
rect 17234 16294 17286 16346
rect 17298 16294 17350 16346
rect 17362 16294 17414 16346
rect 17426 16294 17478 16346
rect 17490 16294 17542 16346
rect 22662 16294 22714 16346
rect 22726 16294 22778 16346
rect 22790 16294 22842 16346
rect 22854 16294 22906 16346
rect 22918 16294 22970 16346
rect 3664 15750 3716 15802
rect 3728 15750 3780 15802
rect 3792 15750 3844 15802
rect 3856 15750 3908 15802
rect 3920 15750 3972 15802
rect 9092 15750 9144 15802
rect 9156 15750 9208 15802
rect 9220 15750 9272 15802
rect 9284 15750 9336 15802
rect 9348 15750 9400 15802
rect 14520 15750 14572 15802
rect 14584 15750 14636 15802
rect 14648 15750 14700 15802
rect 14712 15750 14764 15802
rect 14776 15750 14828 15802
rect 19948 15750 20000 15802
rect 20012 15750 20064 15802
rect 20076 15750 20128 15802
rect 20140 15750 20192 15802
rect 20204 15750 20256 15802
rect 6378 15206 6430 15258
rect 6442 15206 6494 15258
rect 6506 15206 6558 15258
rect 6570 15206 6622 15258
rect 6634 15206 6686 15258
rect 11806 15206 11858 15258
rect 11870 15206 11922 15258
rect 11934 15206 11986 15258
rect 11998 15206 12050 15258
rect 12062 15206 12114 15258
rect 17234 15206 17286 15258
rect 17298 15206 17350 15258
rect 17362 15206 17414 15258
rect 17426 15206 17478 15258
rect 17490 15206 17542 15258
rect 22662 15206 22714 15258
rect 22726 15206 22778 15258
rect 22790 15206 22842 15258
rect 22854 15206 22906 15258
rect 22918 15206 22970 15258
rect 3664 14662 3716 14714
rect 3728 14662 3780 14714
rect 3792 14662 3844 14714
rect 3856 14662 3908 14714
rect 3920 14662 3972 14714
rect 9092 14662 9144 14714
rect 9156 14662 9208 14714
rect 9220 14662 9272 14714
rect 9284 14662 9336 14714
rect 9348 14662 9400 14714
rect 14520 14662 14572 14714
rect 14584 14662 14636 14714
rect 14648 14662 14700 14714
rect 14712 14662 14764 14714
rect 14776 14662 14828 14714
rect 19948 14662 20000 14714
rect 20012 14662 20064 14714
rect 20076 14662 20128 14714
rect 20140 14662 20192 14714
rect 20204 14662 20256 14714
rect 6378 14118 6430 14170
rect 6442 14118 6494 14170
rect 6506 14118 6558 14170
rect 6570 14118 6622 14170
rect 6634 14118 6686 14170
rect 11806 14118 11858 14170
rect 11870 14118 11922 14170
rect 11934 14118 11986 14170
rect 11998 14118 12050 14170
rect 12062 14118 12114 14170
rect 17234 14118 17286 14170
rect 17298 14118 17350 14170
rect 17362 14118 17414 14170
rect 17426 14118 17478 14170
rect 17490 14118 17542 14170
rect 22662 14118 22714 14170
rect 22726 14118 22778 14170
rect 22790 14118 22842 14170
rect 22854 14118 22906 14170
rect 22918 14118 22970 14170
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 17040 13880 17092 13932
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 3664 13574 3716 13626
rect 3728 13574 3780 13626
rect 3792 13574 3844 13626
rect 3856 13574 3908 13626
rect 3920 13574 3972 13626
rect 9092 13574 9144 13626
rect 9156 13574 9208 13626
rect 9220 13574 9272 13626
rect 9284 13574 9336 13626
rect 9348 13574 9400 13626
rect 14520 13574 14572 13626
rect 14584 13574 14636 13626
rect 14648 13574 14700 13626
rect 14712 13574 14764 13626
rect 14776 13574 14828 13626
rect 19948 13574 20000 13626
rect 20012 13574 20064 13626
rect 20076 13574 20128 13626
rect 20140 13574 20192 13626
rect 20204 13574 20256 13626
rect 16212 13268 16264 13320
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 17960 13268 18012 13320
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 8392 13132 8444 13184
rect 17684 13175 17736 13184
rect 17684 13141 17693 13175
rect 17693 13141 17727 13175
rect 17727 13141 17736 13175
rect 17684 13132 17736 13141
rect 19432 13132 19484 13184
rect 6378 13030 6430 13082
rect 6442 13030 6494 13082
rect 6506 13030 6558 13082
rect 6570 13030 6622 13082
rect 6634 13030 6686 13082
rect 11806 13030 11858 13082
rect 11870 13030 11922 13082
rect 11934 13030 11986 13082
rect 11998 13030 12050 13082
rect 12062 13030 12114 13082
rect 17234 13030 17286 13082
rect 17298 13030 17350 13082
rect 17362 13030 17414 13082
rect 17426 13030 17478 13082
rect 17490 13030 17542 13082
rect 22662 13030 22714 13082
rect 22726 13030 22778 13082
rect 22790 13030 22842 13082
rect 22854 13030 22906 13082
rect 22918 13030 22970 13082
rect 16212 12971 16264 12980
rect 16212 12937 16221 12971
rect 16221 12937 16255 12971
rect 16255 12937 16264 12971
rect 16212 12928 16264 12937
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 17960 12792 18012 12844
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 19064 12835 19116 12844
rect 18788 12792 18840 12801
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 20444 12792 20496 12844
rect 17868 12724 17920 12776
rect 18144 12631 18196 12640
rect 18144 12597 18153 12631
rect 18153 12597 18187 12631
rect 18187 12597 18196 12631
rect 18144 12588 18196 12597
rect 18696 12588 18748 12640
rect 18972 12588 19024 12640
rect 3664 12486 3716 12538
rect 3728 12486 3780 12538
rect 3792 12486 3844 12538
rect 3856 12486 3908 12538
rect 3920 12486 3972 12538
rect 9092 12486 9144 12538
rect 9156 12486 9208 12538
rect 9220 12486 9272 12538
rect 9284 12486 9336 12538
rect 9348 12486 9400 12538
rect 14520 12486 14572 12538
rect 14584 12486 14636 12538
rect 14648 12486 14700 12538
rect 14712 12486 14764 12538
rect 14776 12486 14828 12538
rect 19948 12486 20000 12538
rect 20012 12486 20064 12538
rect 20076 12486 20128 12538
rect 20140 12486 20192 12538
rect 20204 12486 20256 12538
rect 16120 12384 16172 12436
rect 18236 12384 18288 12436
rect 18696 12384 18748 12436
rect 20444 12427 20496 12436
rect 20444 12393 20453 12427
rect 20453 12393 20487 12427
rect 20487 12393 20496 12427
rect 20444 12384 20496 12393
rect 18880 12316 18932 12368
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 16028 12180 16080 12232
rect 16948 12180 17000 12232
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 16856 12112 16908 12164
rect 18788 12112 18840 12164
rect 18972 12112 19024 12164
rect 6184 12044 6236 12096
rect 18052 12044 18104 12096
rect 6378 11942 6430 11994
rect 6442 11942 6494 11994
rect 6506 11942 6558 11994
rect 6570 11942 6622 11994
rect 6634 11942 6686 11994
rect 11806 11942 11858 11994
rect 11870 11942 11922 11994
rect 11934 11942 11986 11994
rect 11998 11942 12050 11994
rect 12062 11942 12114 11994
rect 17234 11942 17286 11994
rect 17298 11942 17350 11994
rect 17362 11942 17414 11994
rect 17426 11942 17478 11994
rect 17490 11942 17542 11994
rect 22662 11942 22714 11994
rect 22726 11942 22778 11994
rect 22790 11942 22842 11994
rect 22854 11942 22906 11994
rect 22918 11942 22970 11994
rect 19064 11840 19116 11892
rect 16948 11772 17000 11824
rect 17592 11704 17644 11756
rect 16948 11679 17000 11688
rect 16948 11645 16957 11679
rect 16957 11645 16991 11679
rect 16991 11645 17000 11679
rect 16948 11636 17000 11645
rect 18880 11679 18932 11688
rect 18880 11645 18889 11679
rect 18889 11645 18923 11679
rect 18923 11645 18932 11679
rect 18880 11636 18932 11645
rect 18972 11568 19024 11620
rect 16856 11500 16908 11552
rect 3664 11398 3716 11450
rect 3728 11398 3780 11450
rect 3792 11398 3844 11450
rect 3856 11398 3908 11450
rect 3920 11398 3972 11450
rect 9092 11398 9144 11450
rect 9156 11398 9208 11450
rect 9220 11398 9272 11450
rect 9284 11398 9336 11450
rect 9348 11398 9400 11450
rect 14520 11398 14572 11450
rect 14584 11398 14636 11450
rect 14648 11398 14700 11450
rect 14712 11398 14764 11450
rect 14776 11398 14828 11450
rect 19948 11398 20000 11450
rect 20012 11398 20064 11450
rect 20076 11398 20128 11450
rect 20140 11398 20192 11450
rect 20204 11398 20256 11450
rect 16948 11296 17000 11348
rect 21548 11228 21600 11280
rect 18236 11092 18288 11144
rect 18696 11092 18748 11144
rect 19248 11024 19300 11076
rect 17868 10999 17920 11008
rect 17868 10965 17877 10999
rect 17877 10965 17911 10999
rect 17911 10965 17920 10999
rect 17868 10956 17920 10965
rect 17960 10956 18012 11008
rect 6378 10854 6430 10906
rect 6442 10854 6494 10906
rect 6506 10854 6558 10906
rect 6570 10854 6622 10906
rect 6634 10854 6686 10906
rect 11806 10854 11858 10906
rect 11870 10854 11922 10906
rect 11934 10854 11986 10906
rect 11998 10854 12050 10906
rect 12062 10854 12114 10906
rect 17234 10854 17286 10906
rect 17298 10854 17350 10906
rect 17362 10854 17414 10906
rect 17426 10854 17478 10906
rect 17490 10854 17542 10906
rect 22662 10854 22714 10906
rect 22726 10854 22778 10906
rect 22790 10854 22842 10906
rect 22854 10854 22906 10906
rect 22918 10854 22970 10906
rect 18880 10752 18932 10804
rect 17592 10659 17644 10668
rect 17592 10625 17601 10659
rect 17601 10625 17635 10659
rect 17635 10625 17644 10659
rect 17868 10659 17920 10668
rect 17592 10616 17644 10625
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 19708 10684 19760 10736
rect 18972 10616 19024 10668
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 21364 10616 21416 10668
rect 21180 10480 21232 10532
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 17224 10412 17276 10464
rect 21272 10412 21324 10464
rect 3664 10310 3716 10362
rect 3728 10310 3780 10362
rect 3792 10310 3844 10362
rect 3856 10310 3908 10362
rect 3920 10310 3972 10362
rect 9092 10310 9144 10362
rect 9156 10310 9208 10362
rect 9220 10310 9272 10362
rect 9284 10310 9336 10362
rect 9348 10310 9400 10362
rect 14520 10310 14572 10362
rect 14584 10310 14636 10362
rect 14648 10310 14700 10362
rect 14712 10310 14764 10362
rect 14776 10310 14828 10362
rect 19948 10310 20000 10362
rect 20012 10310 20064 10362
rect 20076 10310 20128 10362
rect 20140 10310 20192 10362
rect 20204 10310 20256 10362
rect 16856 10140 16908 10192
rect 11704 10072 11756 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 18880 10208 18932 10260
rect 19800 10208 19852 10260
rect 18052 10115 18104 10124
rect 18052 10081 18086 10115
rect 18086 10081 18104 10115
rect 18052 10072 18104 10081
rect 18972 10072 19024 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 21548 10115 21600 10124
rect 21548 10081 21557 10115
rect 21557 10081 21591 10115
rect 21591 10081 21600 10115
rect 21548 10072 21600 10081
rect 19432 10047 19484 10056
rect 2504 9868 2556 9920
rect 16856 9868 16908 9920
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 17684 9868 17736 9920
rect 19984 9936 20036 9988
rect 18880 9911 18932 9920
rect 18880 9877 18889 9911
rect 18889 9877 18923 9911
rect 18923 9877 18932 9911
rect 18880 9868 18932 9877
rect 6378 9766 6430 9818
rect 6442 9766 6494 9818
rect 6506 9766 6558 9818
rect 6570 9766 6622 9818
rect 6634 9766 6686 9818
rect 11806 9766 11858 9818
rect 11870 9766 11922 9818
rect 11934 9766 11986 9818
rect 11998 9766 12050 9818
rect 12062 9766 12114 9818
rect 17234 9766 17286 9818
rect 17298 9766 17350 9818
rect 17362 9766 17414 9818
rect 17426 9766 17478 9818
rect 17490 9766 17542 9818
rect 22662 9766 22714 9818
rect 22726 9766 22778 9818
rect 22790 9766 22842 9818
rect 22854 9766 22906 9818
rect 22918 9766 22970 9818
rect 18052 9664 18104 9716
rect 18604 9664 18656 9716
rect 19432 9707 19484 9716
rect 19432 9673 19441 9707
rect 19441 9673 19475 9707
rect 19475 9673 19484 9707
rect 19432 9664 19484 9673
rect 19984 9707 20036 9716
rect 19984 9673 19993 9707
rect 19993 9673 20027 9707
rect 20027 9673 20036 9707
rect 19984 9664 20036 9673
rect 18696 9571 18748 9580
rect 18696 9537 18705 9571
rect 18705 9537 18739 9571
rect 18739 9537 18748 9571
rect 18696 9528 18748 9537
rect 19248 9528 19300 9580
rect 21364 9596 21416 9648
rect 21180 9571 21232 9580
rect 21180 9537 21189 9571
rect 21189 9537 21223 9571
rect 21223 9537 21232 9571
rect 21180 9528 21232 9537
rect 20352 9460 20404 9512
rect 3664 9222 3716 9274
rect 3728 9222 3780 9274
rect 3792 9222 3844 9274
rect 3856 9222 3908 9274
rect 3920 9222 3972 9274
rect 9092 9222 9144 9274
rect 9156 9222 9208 9274
rect 9220 9222 9272 9274
rect 9284 9222 9336 9274
rect 9348 9222 9400 9274
rect 14520 9222 14572 9274
rect 14584 9222 14636 9274
rect 14648 9222 14700 9274
rect 14712 9222 14764 9274
rect 14776 9222 14828 9274
rect 19948 9222 20000 9274
rect 20012 9222 20064 9274
rect 20076 9222 20128 9274
rect 20140 9222 20192 9274
rect 20204 9222 20256 9274
rect 20536 8780 20588 8832
rect 21640 8780 21692 8832
rect 6378 8678 6430 8730
rect 6442 8678 6494 8730
rect 6506 8678 6558 8730
rect 6570 8678 6622 8730
rect 6634 8678 6686 8730
rect 11806 8678 11858 8730
rect 11870 8678 11922 8730
rect 11934 8678 11986 8730
rect 11998 8678 12050 8730
rect 12062 8678 12114 8730
rect 17234 8678 17286 8730
rect 17298 8678 17350 8730
rect 17362 8678 17414 8730
rect 17426 8678 17478 8730
rect 17490 8678 17542 8730
rect 22662 8678 22714 8730
rect 22726 8678 22778 8730
rect 22790 8678 22842 8730
rect 22854 8678 22906 8730
rect 22918 8678 22970 8730
rect 21640 8576 21692 8628
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 20352 8440 20404 8492
rect 20536 8415 20588 8424
rect 20536 8381 20545 8415
rect 20545 8381 20579 8415
rect 20579 8381 20588 8415
rect 20536 8372 20588 8381
rect 18604 8304 18656 8356
rect 20996 8347 21048 8356
rect 18880 8279 18932 8288
rect 18880 8245 18889 8279
rect 18889 8245 18923 8279
rect 18923 8245 18932 8279
rect 18880 8236 18932 8245
rect 20444 8279 20496 8288
rect 20444 8245 20453 8279
rect 20453 8245 20487 8279
rect 20487 8245 20496 8279
rect 20444 8236 20496 8245
rect 20996 8313 21005 8347
rect 21005 8313 21039 8347
rect 21039 8313 21048 8347
rect 20996 8304 21048 8313
rect 21548 8236 21600 8288
rect 3664 8134 3716 8186
rect 3728 8134 3780 8186
rect 3792 8134 3844 8186
rect 3856 8134 3908 8186
rect 3920 8134 3972 8186
rect 9092 8134 9144 8186
rect 9156 8134 9208 8186
rect 9220 8134 9272 8186
rect 9284 8134 9336 8186
rect 9348 8134 9400 8186
rect 14520 8134 14572 8186
rect 14584 8134 14636 8186
rect 14648 8134 14700 8186
rect 14712 8134 14764 8186
rect 14776 8134 14828 8186
rect 19948 8134 20000 8186
rect 20012 8134 20064 8186
rect 20076 8134 20128 8186
rect 20140 8134 20192 8186
rect 20204 8134 20256 8186
rect 18144 7896 18196 7948
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 18696 7760 18748 7812
rect 19156 7760 19208 7812
rect 18512 7692 18564 7744
rect 6378 7590 6430 7642
rect 6442 7590 6494 7642
rect 6506 7590 6558 7642
rect 6570 7590 6622 7642
rect 6634 7590 6686 7642
rect 11806 7590 11858 7642
rect 11870 7590 11922 7642
rect 11934 7590 11986 7642
rect 11998 7590 12050 7642
rect 12062 7590 12114 7642
rect 17234 7590 17286 7642
rect 17298 7590 17350 7642
rect 17362 7590 17414 7642
rect 17426 7590 17478 7642
rect 17490 7590 17542 7642
rect 22662 7590 22714 7642
rect 22726 7590 22778 7642
rect 22790 7590 22842 7642
rect 22854 7590 22906 7642
rect 22918 7590 22970 7642
rect 19248 7488 19300 7540
rect 18052 7420 18104 7472
rect 20536 7420 20588 7472
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 18420 7327 18472 7336
rect 18420 7293 18429 7327
rect 18429 7293 18463 7327
rect 18463 7293 18472 7327
rect 18420 7284 18472 7293
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 9092 7046 9144 7098
rect 9156 7046 9208 7098
rect 9220 7046 9272 7098
rect 9284 7046 9336 7098
rect 9348 7046 9400 7098
rect 14520 7046 14572 7098
rect 14584 7046 14636 7098
rect 14648 7046 14700 7098
rect 14712 7046 14764 7098
rect 14776 7046 14828 7098
rect 19948 7046 20000 7098
rect 20012 7046 20064 7098
rect 20076 7046 20128 7098
rect 20140 7046 20192 7098
rect 20204 7046 20256 7098
rect 6378 6502 6430 6554
rect 6442 6502 6494 6554
rect 6506 6502 6558 6554
rect 6570 6502 6622 6554
rect 6634 6502 6686 6554
rect 11806 6502 11858 6554
rect 11870 6502 11922 6554
rect 11934 6502 11986 6554
rect 11998 6502 12050 6554
rect 12062 6502 12114 6554
rect 17234 6502 17286 6554
rect 17298 6502 17350 6554
rect 17362 6502 17414 6554
rect 17426 6502 17478 6554
rect 17490 6502 17542 6554
rect 22662 6502 22714 6554
rect 22726 6502 22778 6554
rect 22790 6502 22842 6554
rect 22854 6502 22906 6554
rect 22918 6502 22970 6554
rect 21180 6400 21232 6452
rect 20444 6332 20496 6384
rect 20444 6060 20496 6112
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 9092 5958 9144 6010
rect 9156 5958 9208 6010
rect 9220 5958 9272 6010
rect 9284 5958 9336 6010
rect 9348 5958 9400 6010
rect 14520 5958 14572 6010
rect 14584 5958 14636 6010
rect 14648 5958 14700 6010
rect 14712 5958 14764 6010
rect 14776 5958 14828 6010
rect 19948 5958 20000 6010
rect 20012 5958 20064 6010
rect 20076 5958 20128 6010
rect 20140 5958 20192 6010
rect 20204 5958 20256 6010
rect 19340 5652 19392 5704
rect 19616 5584 19668 5636
rect 18236 5516 18288 5568
rect 6378 5414 6430 5466
rect 6442 5414 6494 5466
rect 6506 5414 6558 5466
rect 6570 5414 6622 5466
rect 6634 5414 6686 5466
rect 11806 5414 11858 5466
rect 11870 5414 11922 5466
rect 11934 5414 11986 5466
rect 11998 5414 12050 5466
rect 12062 5414 12114 5466
rect 17234 5414 17286 5466
rect 17298 5414 17350 5466
rect 17362 5414 17414 5466
rect 17426 5414 17478 5466
rect 17490 5414 17542 5466
rect 22662 5414 22714 5466
rect 22726 5414 22778 5466
rect 22790 5414 22842 5466
rect 22854 5414 22906 5466
rect 22918 5414 22970 5466
rect 20444 5312 20496 5364
rect 20812 5244 20864 5296
rect 19340 5176 19392 5228
rect 19340 4972 19392 5024
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 9092 4870 9144 4922
rect 9156 4870 9208 4922
rect 9220 4870 9272 4922
rect 9284 4870 9336 4922
rect 9348 4870 9400 4922
rect 14520 4870 14572 4922
rect 14584 4870 14636 4922
rect 14648 4870 14700 4922
rect 14712 4870 14764 4922
rect 14776 4870 14828 4922
rect 19948 4870 20000 4922
rect 20012 4870 20064 4922
rect 20076 4870 20128 4922
rect 20140 4870 20192 4922
rect 20204 4870 20256 4922
rect 19616 4768 19668 4820
rect 15660 4700 15712 4752
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 18512 4539 18564 4548
rect 18512 4505 18521 4539
rect 18521 4505 18555 4539
rect 18555 4505 18564 4539
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 20536 4768 20588 4820
rect 19616 4564 19668 4573
rect 22100 4564 22152 4616
rect 18512 4496 18564 4505
rect 22008 4496 22060 4548
rect 22192 4471 22244 4480
rect 22192 4437 22201 4471
rect 22201 4437 22235 4471
rect 22235 4437 22244 4471
rect 22192 4428 22244 4437
rect 6378 4326 6430 4378
rect 6442 4326 6494 4378
rect 6506 4326 6558 4378
rect 6570 4326 6622 4378
rect 6634 4326 6686 4378
rect 11806 4326 11858 4378
rect 11870 4326 11922 4378
rect 11934 4326 11986 4378
rect 11998 4326 12050 4378
rect 12062 4326 12114 4378
rect 17234 4326 17286 4378
rect 17298 4326 17350 4378
rect 17362 4326 17414 4378
rect 17426 4326 17478 4378
rect 17490 4326 17542 4378
rect 22662 4326 22714 4378
rect 22726 4326 22778 4378
rect 22790 4326 22842 4378
rect 22854 4326 22906 4378
rect 22918 4326 22970 4378
rect 19340 4131 19392 4140
rect 19340 4097 19349 4131
rect 19349 4097 19383 4131
rect 19383 4097 19392 4131
rect 19340 4088 19392 4097
rect 19524 4088 19576 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 9092 3782 9144 3834
rect 9156 3782 9208 3834
rect 9220 3782 9272 3834
rect 9284 3782 9336 3834
rect 9348 3782 9400 3834
rect 14520 3782 14572 3834
rect 14584 3782 14636 3834
rect 14648 3782 14700 3834
rect 14712 3782 14764 3834
rect 14776 3782 14828 3834
rect 19948 3782 20000 3834
rect 20012 3782 20064 3834
rect 20076 3782 20128 3834
rect 20140 3782 20192 3834
rect 20204 3782 20256 3834
rect 19524 3680 19576 3732
rect 20812 3723 20864 3732
rect 20812 3689 20821 3723
rect 20821 3689 20855 3723
rect 20855 3689 20864 3723
rect 20812 3680 20864 3689
rect 21364 3544 21416 3596
rect 19616 3476 19668 3528
rect 21824 3408 21876 3460
rect 22192 3408 22244 3460
rect 12992 3340 13044 3392
rect 14372 3340 14424 3392
rect 6378 3238 6430 3290
rect 6442 3238 6494 3290
rect 6506 3238 6558 3290
rect 6570 3238 6622 3290
rect 6634 3238 6686 3290
rect 11806 3238 11858 3290
rect 11870 3238 11922 3290
rect 11934 3238 11986 3290
rect 11998 3238 12050 3290
rect 12062 3238 12114 3290
rect 17234 3238 17286 3290
rect 17298 3238 17350 3290
rect 17362 3238 17414 3290
rect 17426 3238 17478 3290
rect 17490 3238 17542 3290
rect 22662 3238 22714 3290
rect 22726 3238 22778 3290
rect 22790 3238 22842 3290
rect 22854 3238 22906 3290
rect 22918 3238 22970 3290
rect 18420 3136 18472 3188
rect 22100 3179 22152 3188
rect 22100 3145 22109 3179
rect 22109 3145 22143 3179
rect 22143 3145 22152 3179
rect 22100 3136 22152 3145
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 14096 3043 14148 3052
rect 12348 2932 12400 2984
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 13360 2796 13412 2848
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 18236 3068 18288 3120
rect 14372 3000 14424 3009
rect 15660 2864 15712 2916
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 17868 2796 17920 2848
rect 19708 2932 19760 2984
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 9092 2694 9144 2746
rect 9156 2694 9208 2746
rect 9220 2694 9272 2746
rect 9284 2694 9336 2746
rect 9348 2694 9400 2746
rect 14520 2694 14572 2746
rect 14584 2694 14636 2746
rect 14648 2694 14700 2746
rect 14712 2694 14764 2746
rect 14776 2694 14828 2746
rect 19948 2694 20000 2746
rect 20012 2694 20064 2746
rect 20076 2694 20128 2746
rect 20140 2694 20192 2746
rect 20204 2694 20256 2746
rect 12348 2592 12400 2644
rect 14096 2592 14148 2644
rect 18880 2592 18932 2644
rect 12992 2524 13044 2576
rect 2044 2388 2096 2440
rect 6000 2388 6052 2440
rect 9956 2388 10008 2440
rect 13912 2388 13964 2440
rect 20812 2388 20864 2440
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 20996 2320 21048 2372
rect 13360 2252 13412 2304
rect 6378 2150 6430 2202
rect 6442 2150 6494 2202
rect 6506 2150 6558 2202
rect 6570 2150 6622 2202
rect 6634 2150 6686 2202
rect 11806 2150 11858 2202
rect 11870 2150 11922 2202
rect 11934 2150 11986 2202
rect 11998 2150 12050 2202
rect 12062 2150 12114 2202
rect 17234 2150 17286 2202
rect 17298 2150 17350 2202
rect 17362 2150 17414 2202
rect 17426 2150 17478 2202
rect 17490 2150 17542 2202
rect 22662 2150 22714 2202
rect 22726 2150 22778 2202
rect 22790 2150 22842 2202
rect 22854 2150 22906 2202
rect 22918 2150 22970 2202
<< metal2 >>
rect 1674 23338 1730 24000
rect 4618 23338 4674 24000
rect 7562 23338 7618 24000
rect 10506 23338 10562 24000
rect 13450 23338 13506 24000
rect 16394 23338 16450 24000
rect 19338 23338 19394 24000
rect 22282 23338 22338 24000
rect 1674 23310 1900 23338
rect 1674 23200 1730 23310
rect 1872 21690 1900 23310
rect 4618 23310 4844 23338
rect 4618 23200 4674 23310
rect 4816 21690 4844 23310
rect 7562 23310 7788 23338
rect 7562 23200 7618 23310
rect 6378 21788 6686 21797
rect 6378 21786 6384 21788
rect 6440 21786 6464 21788
rect 6520 21786 6544 21788
rect 6600 21786 6624 21788
rect 6680 21786 6686 21788
rect 6440 21734 6442 21786
rect 6622 21734 6624 21786
rect 6378 21732 6384 21734
rect 6440 21732 6464 21734
rect 6520 21732 6544 21734
rect 6600 21732 6624 21734
rect 6680 21732 6686 21734
rect 6378 21723 6686 21732
rect 7760 21690 7788 23310
rect 10506 23310 10732 23338
rect 10506 23200 10562 23310
rect 10704 21690 10732 23310
rect 13450 23310 13768 23338
rect 13450 23200 13506 23310
rect 11806 21788 12114 21797
rect 11806 21786 11812 21788
rect 11868 21786 11892 21788
rect 11948 21786 11972 21788
rect 12028 21786 12052 21788
rect 12108 21786 12114 21788
rect 11868 21734 11870 21786
rect 12050 21734 12052 21786
rect 11806 21732 11812 21734
rect 11868 21732 11892 21734
rect 11948 21732 11972 21734
rect 12028 21732 12052 21734
rect 12108 21732 12114 21734
rect 11806 21723 12114 21732
rect 1860 21684 1912 21690
rect 1860 21626 1912 21632
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 10692 21684 10744 21690
rect 13740 21672 13768 23310
rect 16394 23310 16528 23338
rect 16394 23200 16450 23310
rect 13820 21684 13872 21690
rect 13740 21644 13820 21672
rect 10692 21626 10744 21632
rect 16500 21672 16528 23310
rect 19338 23310 19564 23338
rect 19338 23200 19394 23310
rect 17234 21788 17542 21797
rect 17234 21786 17240 21788
rect 17296 21786 17320 21788
rect 17376 21786 17400 21788
rect 17456 21786 17480 21788
rect 17536 21786 17542 21788
rect 17296 21734 17298 21786
rect 17478 21734 17480 21786
rect 17234 21732 17240 21734
rect 17296 21732 17320 21734
rect 17376 21732 17400 21734
rect 17456 21732 17480 21734
rect 17536 21732 17542 21734
rect 17234 21723 17542 21732
rect 19536 21690 19564 23310
rect 22204 23310 22338 23338
rect 22204 21690 22232 23310
rect 22282 23200 22338 23310
rect 22662 21788 22970 21797
rect 22662 21786 22668 21788
rect 22724 21786 22748 21788
rect 22804 21786 22828 21788
rect 22884 21786 22908 21788
rect 22964 21786 22970 21788
rect 22724 21734 22726 21786
rect 22906 21734 22908 21786
rect 22662 21732 22668 21734
rect 22724 21732 22748 21734
rect 22804 21732 22828 21734
rect 22884 21732 22908 21734
rect 22964 21732 22970 21734
rect 22662 21723 22970 21732
rect 16580 21684 16632 21690
rect 16500 21644 16580 21672
rect 13820 21626 13872 21632
rect 16580 21626 16632 21632
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 2516 21350 2544 21490
rect 8404 21350 8432 21490
rect 11716 21350 11744 21490
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 2516 9926 2544 21286
rect 3664 21244 3972 21253
rect 3664 21242 3670 21244
rect 3726 21242 3750 21244
rect 3806 21242 3830 21244
rect 3886 21242 3910 21244
rect 3966 21242 3972 21244
rect 3726 21190 3728 21242
rect 3908 21190 3910 21242
rect 3664 21188 3670 21190
rect 3726 21188 3750 21190
rect 3806 21188 3830 21190
rect 3886 21188 3910 21190
rect 3966 21188 3972 21190
rect 3664 21179 3972 21188
rect 3664 20156 3972 20165
rect 3664 20154 3670 20156
rect 3726 20154 3750 20156
rect 3806 20154 3830 20156
rect 3886 20154 3910 20156
rect 3966 20154 3972 20156
rect 3726 20102 3728 20154
rect 3908 20102 3910 20154
rect 3664 20100 3670 20102
rect 3726 20100 3750 20102
rect 3806 20100 3830 20102
rect 3886 20100 3910 20102
rect 3966 20100 3972 20102
rect 3664 20091 3972 20100
rect 3664 19068 3972 19077
rect 3664 19066 3670 19068
rect 3726 19066 3750 19068
rect 3806 19066 3830 19068
rect 3886 19066 3910 19068
rect 3966 19066 3972 19068
rect 3726 19014 3728 19066
rect 3908 19014 3910 19066
rect 3664 19012 3670 19014
rect 3726 19012 3750 19014
rect 3806 19012 3830 19014
rect 3886 19012 3910 19014
rect 3966 19012 3972 19014
rect 3664 19003 3972 19012
rect 3664 17980 3972 17989
rect 3664 17978 3670 17980
rect 3726 17978 3750 17980
rect 3806 17978 3830 17980
rect 3886 17978 3910 17980
rect 3966 17978 3972 17980
rect 3726 17926 3728 17978
rect 3908 17926 3910 17978
rect 3664 17924 3670 17926
rect 3726 17924 3750 17926
rect 3806 17924 3830 17926
rect 3886 17924 3910 17926
rect 3966 17924 3972 17926
rect 3664 17915 3972 17924
rect 3664 16892 3972 16901
rect 3664 16890 3670 16892
rect 3726 16890 3750 16892
rect 3806 16890 3830 16892
rect 3886 16890 3910 16892
rect 3966 16890 3972 16892
rect 3726 16838 3728 16890
rect 3908 16838 3910 16890
rect 3664 16836 3670 16838
rect 3726 16836 3750 16838
rect 3806 16836 3830 16838
rect 3886 16836 3910 16838
rect 3966 16836 3972 16838
rect 3664 16827 3972 16836
rect 3664 15804 3972 15813
rect 3664 15802 3670 15804
rect 3726 15802 3750 15804
rect 3806 15802 3830 15804
rect 3886 15802 3910 15804
rect 3966 15802 3972 15804
rect 3726 15750 3728 15802
rect 3908 15750 3910 15802
rect 3664 15748 3670 15750
rect 3726 15748 3750 15750
rect 3806 15748 3830 15750
rect 3886 15748 3910 15750
rect 3966 15748 3972 15750
rect 3664 15739 3972 15748
rect 3664 14716 3972 14725
rect 3664 14714 3670 14716
rect 3726 14714 3750 14716
rect 3806 14714 3830 14716
rect 3886 14714 3910 14716
rect 3966 14714 3972 14716
rect 3726 14662 3728 14714
rect 3908 14662 3910 14714
rect 3664 14660 3670 14662
rect 3726 14660 3750 14662
rect 3806 14660 3830 14662
rect 3886 14660 3910 14662
rect 3966 14660 3972 14662
rect 3664 14651 3972 14660
rect 3664 13628 3972 13637
rect 3664 13626 3670 13628
rect 3726 13626 3750 13628
rect 3806 13626 3830 13628
rect 3886 13626 3910 13628
rect 3966 13626 3972 13628
rect 3726 13574 3728 13626
rect 3908 13574 3910 13626
rect 3664 13572 3670 13574
rect 3726 13572 3750 13574
rect 3806 13572 3830 13574
rect 3886 13572 3910 13574
rect 3966 13572 3972 13574
rect 3664 13563 3972 13572
rect 3664 12540 3972 12549
rect 3664 12538 3670 12540
rect 3726 12538 3750 12540
rect 3806 12538 3830 12540
rect 3886 12538 3910 12540
rect 3966 12538 3972 12540
rect 3726 12486 3728 12538
rect 3908 12486 3910 12538
rect 3664 12484 3670 12486
rect 3726 12484 3750 12486
rect 3806 12484 3830 12486
rect 3886 12484 3910 12486
rect 3966 12484 3972 12486
rect 3664 12475 3972 12484
rect 6196 12102 6224 21286
rect 6378 20700 6686 20709
rect 6378 20698 6384 20700
rect 6440 20698 6464 20700
rect 6520 20698 6544 20700
rect 6600 20698 6624 20700
rect 6680 20698 6686 20700
rect 6440 20646 6442 20698
rect 6622 20646 6624 20698
rect 6378 20644 6384 20646
rect 6440 20644 6464 20646
rect 6520 20644 6544 20646
rect 6600 20644 6624 20646
rect 6680 20644 6686 20646
rect 6378 20635 6686 20644
rect 6378 19612 6686 19621
rect 6378 19610 6384 19612
rect 6440 19610 6464 19612
rect 6520 19610 6544 19612
rect 6600 19610 6624 19612
rect 6680 19610 6686 19612
rect 6440 19558 6442 19610
rect 6622 19558 6624 19610
rect 6378 19556 6384 19558
rect 6440 19556 6464 19558
rect 6520 19556 6544 19558
rect 6600 19556 6624 19558
rect 6680 19556 6686 19558
rect 6378 19547 6686 19556
rect 6378 18524 6686 18533
rect 6378 18522 6384 18524
rect 6440 18522 6464 18524
rect 6520 18522 6544 18524
rect 6600 18522 6624 18524
rect 6680 18522 6686 18524
rect 6440 18470 6442 18522
rect 6622 18470 6624 18522
rect 6378 18468 6384 18470
rect 6440 18468 6464 18470
rect 6520 18468 6544 18470
rect 6600 18468 6624 18470
rect 6680 18468 6686 18470
rect 6378 18459 6686 18468
rect 6378 17436 6686 17445
rect 6378 17434 6384 17436
rect 6440 17434 6464 17436
rect 6520 17434 6544 17436
rect 6600 17434 6624 17436
rect 6680 17434 6686 17436
rect 6440 17382 6442 17434
rect 6622 17382 6624 17434
rect 6378 17380 6384 17382
rect 6440 17380 6464 17382
rect 6520 17380 6544 17382
rect 6600 17380 6624 17382
rect 6680 17380 6686 17382
rect 6378 17371 6686 17380
rect 6378 16348 6686 16357
rect 6378 16346 6384 16348
rect 6440 16346 6464 16348
rect 6520 16346 6544 16348
rect 6600 16346 6624 16348
rect 6680 16346 6686 16348
rect 6440 16294 6442 16346
rect 6622 16294 6624 16346
rect 6378 16292 6384 16294
rect 6440 16292 6464 16294
rect 6520 16292 6544 16294
rect 6600 16292 6624 16294
rect 6680 16292 6686 16294
rect 6378 16283 6686 16292
rect 6378 15260 6686 15269
rect 6378 15258 6384 15260
rect 6440 15258 6464 15260
rect 6520 15258 6544 15260
rect 6600 15258 6624 15260
rect 6680 15258 6686 15260
rect 6440 15206 6442 15258
rect 6622 15206 6624 15258
rect 6378 15204 6384 15206
rect 6440 15204 6464 15206
rect 6520 15204 6544 15206
rect 6600 15204 6624 15206
rect 6680 15204 6686 15206
rect 6378 15195 6686 15204
rect 6378 14172 6686 14181
rect 6378 14170 6384 14172
rect 6440 14170 6464 14172
rect 6520 14170 6544 14172
rect 6600 14170 6624 14172
rect 6680 14170 6686 14172
rect 6440 14118 6442 14170
rect 6622 14118 6624 14170
rect 6378 14116 6384 14118
rect 6440 14116 6464 14118
rect 6520 14116 6544 14118
rect 6600 14116 6624 14118
rect 6680 14116 6686 14118
rect 6378 14107 6686 14116
rect 8404 13190 8432 21286
rect 9092 21244 9400 21253
rect 9092 21242 9098 21244
rect 9154 21242 9178 21244
rect 9234 21242 9258 21244
rect 9314 21242 9338 21244
rect 9394 21242 9400 21244
rect 9154 21190 9156 21242
rect 9336 21190 9338 21242
rect 9092 21188 9098 21190
rect 9154 21188 9178 21190
rect 9234 21188 9258 21190
rect 9314 21188 9338 21190
rect 9394 21188 9400 21190
rect 9092 21179 9400 21188
rect 9092 20156 9400 20165
rect 9092 20154 9098 20156
rect 9154 20154 9178 20156
rect 9234 20154 9258 20156
rect 9314 20154 9338 20156
rect 9394 20154 9400 20156
rect 9154 20102 9156 20154
rect 9336 20102 9338 20154
rect 9092 20100 9098 20102
rect 9154 20100 9178 20102
rect 9234 20100 9258 20102
rect 9314 20100 9338 20102
rect 9394 20100 9400 20102
rect 9092 20091 9400 20100
rect 9092 19068 9400 19077
rect 9092 19066 9098 19068
rect 9154 19066 9178 19068
rect 9234 19066 9258 19068
rect 9314 19066 9338 19068
rect 9394 19066 9400 19068
rect 9154 19014 9156 19066
rect 9336 19014 9338 19066
rect 9092 19012 9098 19014
rect 9154 19012 9178 19014
rect 9234 19012 9258 19014
rect 9314 19012 9338 19014
rect 9394 19012 9400 19014
rect 9092 19003 9400 19012
rect 9092 17980 9400 17989
rect 9092 17978 9098 17980
rect 9154 17978 9178 17980
rect 9234 17978 9258 17980
rect 9314 17978 9338 17980
rect 9394 17978 9400 17980
rect 9154 17926 9156 17978
rect 9336 17926 9338 17978
rect 9092 17924 9098 17926
rect 9154 17924 9178 17926
rect 9234 17924 9258 17926
rect 9314 17924 9338 17926
rect 9394 17924 9400 17926
rect 9092 17915 9400 17924
rect 9092 16892 9400 16901
rect 9092 16890 9098 16892
rect 9154 16890 9178 16892
rect 9234 16890 9258 16892
rect 9314 16890 9338 16892
rect 9394 16890 9400 16892
rect 9154 16838 9156 16890
rect 9336 16838 9338 16890
rect 9092 16836 9098 16838
rect 9154 16836 9178 16838
rect 9234 16836 9258 16838
rect 9314 16836 9338 16838
rect 9394 16836 9400 16838
rect 9092 16827 9400 16836
rect 9092 15804 9400 15813
rect 9092 15802 9098 15804
rect 9154 15802 9178 15804
rect 9234 15802 9258 15804
rect 9314 15802 9338 15804
rect 9394 15802 9400 15804
rect 9154 15750 9156 15802
rect 9336 15750 9338 15802
rect 9092 15748 9098 15750
rect 9154 15748 9178 15750
rect 9234 15748 9258 15750
rect 9314 15748 9338 15750
rect 9394 15748 9400 15750
rect 9092 15739 9400 15748
rect 9092 14716 9400 14725
rect 9092 14714 9098 14716
rect 9154 14714 9178 14716
rect 9234 14714 9258 14716
rect 9314 14714 9338 14716
rect 9394 14714 9400 14716
rect 9154 14662 9156 14714
rect 9336 14662 9338 14714
rect 9092 14660 9098 14662
rect 9154 14660 9178 14662
rect 9234 14660 9258 14662
rect 9314 14660 9338 14662
rect 9394 14660 9400 14662
rect 9092 14651 9400 14660
rect 9092 13628 9400 13637
rect 9092 13626 9098 13628
rect 9154 13626 9178 13628
rect 9234 13626 9258 13628
rect 9314 13626 9338 13628
rect 9394 13626 9400 13628
rect 9154 13574 9156 13626
rect 9336 13574 9338 13626
rect 9092 13572 9098 13574
rect 9154 13572 9178 13574
rect 9234 13572 9258 13574
rect 9314 13572 9338 13574
rect 9394 13572 9400 13574
rect 9092 13563 9400 13572
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 6378 13084 6686 13093
rect 6378 13082 6384 13084
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6680 13082 6686 13084
rect 6440 13030 6442 13082
rect 6622 13030 6624 13082
rect 6378 13028 6384 13030
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6680 13028 6686 13030
rect 6378 13019 6686 13028
rect 9092 12540 9400 12549
rect 9092 12538 9098 12540
rect 9154 12538 9178 12540
rect 9234 12538 9258 12540
rect 9314 12538 9338 12540
rect 9394 12538 9400 12540
rect 9154 12486 9156 12538
rect 9336 12486 9338 12538
rect 9092 12484 9098 12486
rect 9154 12484 9178 12486
rect 9234 12484 9258 12486
rect 9314 12484 9338 12486
rect 9394 12484 9400 12486
rect 9092 12475 9400 12484
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6378 11996 6686 12005
rect 6378 11994 6384 11996
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6680 11994 6686 11996
rect 6440 11942 6442 11994
rect 6622 11942 6624 11994
rect 6378 11940 6384 11942
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6680 11940 6686 11942
rect 6378 11931 6686 11940
rect 3664 11452 3972 11461
rect 3664 11450 3670 11452
rect 3726 11450 3750 11452
rect 3806 11450 3830 11452
rect 3886 11450 3910 11452
rect 3966 11450 3972 11452
rect 3726 11398 3728 11450
rect 3908 11398 3910 11450
rect 3664 11396 3670 11398
rect 3726 11396 3750 11398
rect 3806 11396 3830 11398
rect 3886 11396 3910 11398
rect 3966 11396 3972 11398
rect 3664 11387 3972 11396
rect 9092 11452 9400 11461
rect 9092 11450 9098 11452
rect 9154 11450 9178 11452
rect 9234 11450 9258 11452
rect 9314 11450 9338 11452
rect 9394 11450 9400 11452
rect 9154 11398 9156 11450
rect 9336 11398 9338 11450
rect 9092 11396 9098 11398
rect 9154 11396 9178 11398
rect 9234 11396 9258 11398
rect 9314 11396 9338 11398
rect 9394 11396 9400 11398
rect 9092 11387 9400 11396
rect 6378 10908 6686 10917
rect 6378 10906 6384 10908
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6680 10906 6686 10908
rect 6440 10854 6442 10906
rect 6622 10854 6624 10906
rect 6378 10852 6384 10854
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6680 10852 6686 10854
rect 6378 10843 6686 10852
rect 3664 10364 3972 10373
rect 3664 10362 3670 10364
rect 3726 10362 3750 10364
rect 3806 10362 3830 10364
rect 3886 10362 3910 10364
rect 3966 10362 3972 10364
rect 3726 10310 3728 10362
rect 3908 10310 3910 10362
rect 3664 10308 3670 10310
rect 3726 10308 3750 10310
rect 3806 10308 3830 10310
rect 3886 10308 3910 10310
rect 3966 10308 3972 10310
rect 3664 10299 3972 10308
rect 9092 10364 9400 10373
rect 9092 10362 9098 10364
rect 9154 10362 9178 10364
rect 9234 10362 9258 10364
rect 9314 10362 9338 10364
rect 9394 10362 9400 10364
rect 9154 10310 9156 10362
rect 9336 10310 9338 10362
rect 9092 10308 9098 10310
rect 9154 10308 9178 10310
rect 9234 10308 9258 10310
rect 9314 10308 9338 10310
rect 9394 10308 9400 10310
rect 9092 10299 9400 10308
rect 11716 10130 11744 21286
rect 14520 21244 14828 21253
rect 14520 21242 14526 21244
rect 14582 21242 14606 21244
rect 14662 21242 14686 21244
rect 14742 21242 14766 21244
rect 14822 21242 14828 21244
rect 14582 21190 14584 21242
rect 14764 21190 14766 21242
rect 14520 21188 14526 21190
rect 14582 21188 14606 21190
rect 14662 21188 14686 21190
rect 14742 21188 14766 21190
rect 14822 21188 14828 21190
rect 14520 21179 14828 21188
rect 11806 20700 12114 20709
rect 11806 20698 11812 20700
rect 11868 20698 11892 20700
rect 11948 20698 11972 20700
rect 12028 20698 12052 20700
rect 12108 20698 12114 20700
rect 11868 20646 11870 20698
rect 12050 20646 12052 20698
rect 11806 20644 11812 20646
rect 11868 20644 11892 20646
rect 11948 20644 11972 20646
rect 12028 20644 12052 20646
rect 12108 20644 12114 20646
rect 11806 20635 12114 20644
rect 17234 20700 17542 20709
rect 17234 20698 17240 20700
rect 17296 20698 17320 20700
rect 17376 20698 17400 20700
rect 17456 20698 17480 20700
rect 17536 20698 17542 20700
rect 17296 20646 17298 20698
rect 17478 20646 17480 20698
rect 17234 20644 17240 20646
rect 17296 20644 17320 20646
rect 17376 20644 17400 20646
rect 17456 20644 17480 20646
rect 17536 20644 17542 20646
rect 17234 20635 17542 20644
rect 14520 20156 14828 20165
rect 14520 20154 14526 20156
rect 14582 20154 14606 20156
rect 14662 20154 14686 20156
rect 14742 20154 14766 20156
rect 14822 20154 14828 20156
rect 14582 20102 14584 20154
rect 14764 20102 14766 20154
rect 14520 20100 14526 20102
rect 14582 20100 14606 20102
rect 14662 20100 14686 20102
rect 14742 20100 14766 20102
rect 14822 20100 14828 20102
rect 14520 20091 14828 20100
rect 11806 19612 12114 19621
rect 11806 19610 11812 19612
rect 11868 19610 11892 19612
rect 11948 19610 11972 19612
rect 12028 19610 12052 19612
rect 12108 19610 12114 19612
rect 11868 19558 11870 19610
rect 12050 19558 12052 19610
rect 11806 19556 11812 19558
rect 11868 19556 11892 19558
rect 11948 19556 11972 19558
rect 12028 19556 12052 19558
rect 12108 19556 12114 19558
rect 11806 19547 12114 19556
rect 17234 19612 17542 19621
rect 17234 19610 17240 19612
rect 17296 19610 17320 19612
rect 17376 19610 17400 19612
rect 17456 19610 17480 19612
rect 17536 19610 17542 19612
rect 17296 19558 17298 19610
rect 17478 19558 17480 19610
rect 17234 19556 17240 19558
rect 17296 19556 17320 19558
rect 17376 19556 17400 19558
rect 17456 19556 17480 19558
rect 17536 19556 17542 19558
rect 17234 19547 17542 19556
rect 14520 19068 14828 19077
rect 14520 19066 14526 19068
rect 14582 19066 14606 19068
rect 14662 19066 14686 19068
rect 14742 19066 14766 19068
rect 14822 19066 14828 19068
rect 14582 19014 14584 19066
rect 14764 19014 14766 19066
rect 14520 19012 14526 19014
rect 14582 19012 14606 19014
rect 14662 19012 14686 19014
rect 14742 19012 14766 19014
rect 14822 19012 14828 19014
rect 14520 19003 14828 19012
rect 11806 18524 12114 18533
rect 11806 18522 11812 18524
rect 11868 18522 11892 18524
rect 11948 18522 11972 18524
rect 12028 18522 12052 18524
rect 12108 18522 12114 18524
rect 11868 18470 11870 18522
rect 12050 18470 12052 18522
rect 11806 18468 11812 18470
rect 11868 18468 11892 18470
rect 11948 18468 11972 18470
rect 12028 18468 12052 18470
rect 12108 18468 12114 18470
rect 11806 18459 12114 18468
rect 17234 18524 17542 18533
rect 17234 18522 17240 18524
rect 17296 18522 17320 18524
rect 17376 18522 17400 18524
rect 17456 18522 17480 18524
rect 17536 18522 17542 18524
rect 17296 18470 17298 18522
rect 17478 18470 17480 18522
rect 17234 18468 17240 18470
rect 17296 18468 17320 18470
rect 17376 18468 17400 18470
rect 17456 18468 17480 18470
rect 17536 18468 17542 18470
rect 17234 18459 17542 18468
rect 14520 17980 14828 17989
rect 14520 17978 14526 17980
rect 14582 17978 14606 17980
rect 14662 17978 14686 17980
rect 14742 17978 14766 17980
rect 14822 17978 14828 17980
rect 14582 17926 14584 17978
rect 14764 17926 14766 17978
rect 14520 17924 14526 17926
rect 14582 17924 14606 17926
rect 14662 17924 14686 17926
rect 14742 17924 14766 17926
rect 14822 17924 14828 17926
rect 14520 17915 14828 17924
rect 11806 17436 12114 17445
rect 11806 17434 11812 17436
rect 11868 17434 11892 17436
rect 11948 17434 11972 17436
rect 12028 17434 12052 17436
rect 12108 17434 12114 17436
rect 11868 17382 11870 17434
rect 12050 17382 12052 17434
rect 11806 17380 11812 17382
rect 11868 17380 11892 17382
rect 11948 17380 11972 17382
rect 12028 17380 12052 17382
rect 12108 17380 12114 17382
rect 11806 17371 12114 17380
rect 17234 17436 17542 17445
rect 17234 17434 17240 17436
rect 17296 17434 17320 17436
rect 17376 17434 17400 17436
rect 17456 17434 17480 17436
rect 17536 17434 17542 17436
rect 17296 17382 17298 17434
rect 17478 17382 17480 17434
rect 17234 17380 17240 17382
rect 17296 17380 17320 17382
rect 17376 17380 17400 17382
rect 17456 17380 17480 17382
rect 17536 17380 17542 17382
rect 17234 17371 17542 17380
rect 14520 16892 14828 16901
rect 14520 16890 14526 16892
rect 14582 16890 14606 16892
rect 14662 16890 14686 16892
rect 14742 16890 14766 16892
rect 14822 16890 14828 16892
rect 14582 16838 14584 16890
rect 14764 16838 14766 16890
rect 14520 16836 14526 16838
rect 14582 16836 14606 16838
rect 14662 16836 14686 16838
rect 14742 16836 14766 16838
rect 14822 16836 14828 16838
rect 14520 16827 14828 16836
rect 11806 16348 12114 16357
rect 11806 16346 11812 16348
rect 11868 16346 11892 16348
rect 11948 16346 11972 16348
rect 12028 16346 12052 16348
rect 12108 16346 12114 16348
rect 11868 16294 11870 16346
rect 12050 16294 12052 16346
rect 11806 16292 11812 16294
rect 11868 16292 11892 16294
rect 11948 16292 11972 16294
rect 12028 16292 12052 16294
rect 12108 16292 12114 16294
rect 11806 16283 12114 16292
rect 17234 16348 17542 16357
rect 17234 16346 17240 16348
rect 17296 16346 17320 16348
rect 17376 16346 17400 16348
rect 17456 16346 17480 16348
rect 17536 16346 17542 16348
rect 17296 16294 17298 16346
rect 17478 16294 17480 16346
rect 17234 16292 17240 16294
rect 17296 16292 17320 16294
rect 17376 16292 17400 16294
rect 17456 16292 17480 16294
rect 17536 16292 17542 16294
rect 17234 16283 17542 16292
rect 14520 15804 14828 15813
rect 14520 15802 14526 15804
rect 14582 15802 14606 15804
rect 14662 15802 14686 15804
rect 14742 15802 14766 15804
rect 14822 15802 14828 15804
rect 14582 15750 14584 15802
rect 14764 15750 14766 15802
rect 14520 15748 14526 15750
rect 14582 15748 14606 15750
rect 14662 15748 14686 15750
rect 14742 15748 14766 15750
rect 14822 15748 14828 15750
rect 14520 15739 14828 15748
rect 11806 15260 12114 15269
rect 11806 15258 11812 15260
rect 11868 15258 11892 15260
rect 11948 15258 11972 15260
rect 12028 15258 12052 15260
rect 12108 15258 12114 15260
rect 11868 15206 11870 15258
rect 12050 15206 12052 15258
rect 11806 15204 11812 15206
rect 11868 15204 11892 15206
rect 11948 15204 11972 15206
rect 12028 15204 12052 15206
rect 12108 15204 12114 15206
rect 11806 15195 12114 15204
rect 17234 15260 17542 15269
rect 17234 15258 17240 15260
rect 17296 15258 17320 15260
rect 17376 15258 17400 15260
rect 17456 15258 17480 15260
rect 17536 15258 17542 15260
rect 17296 15206 17298 15258
rect 17478 15206 17480 15258
rect 17234 15204 17240 15206
rect 17296 15204 17320 15206
rect 17376 15204 17400 15206
rect 17456 15204 17480 15206
rect 17536 15204 17542 15206
rect 17234 15195 17542 15204
rect 14520 14716 14828 14725
rect 14520 14714 14526 14716
rect 14582 14714 14606 14716
rect 14662 14714 14686 14716
rect 14742 14714 14766 14716
rect 14822 14714 14828 14716
rect 14582 14662 14584 14714
rect 14764 14662 14766 14714
rect 14520 14660 14526 14662
rect 14582 14660 14606 14662
rect 14662 14660 14686 14662
rect 14742 14660 14766 14662
rect 14822 14660 14828 14662
rect 14520 14651 14828 14660
rect 11806 14172 12114 14181
rect 11806 14170 11812 14172
rect 11868 14170 11892 14172
rect 11948 14170 11972 14172
rect 12028 14170 12052 14172
rect 12108 14170 12114 14172
rect 11868 14118 11870 14170
rect 12050 14118 12052 14170
rect 11806 14116 11812 14118
rect 11868 14116 11892 14118
rect 11948 14116 11972 14118
rect 12028 14116 12052 14118
rect 12108 14116 12114 14118
rect 11806 14107 12114 14116
rect 17234 14172 17542 14181
rect 17234 14170 17240 14172
rect 17296 14170 17320 14172
rect 17376 14170 17400 14172
rect 17456 14170 17480 14172
rect 17536 14170 17542 14172
rect 17296 14118 17298 14170
rect 17478 14118 17480 14170
rect 17234 14116 17240 14118
rect 17296 14116 17320 14118
rect 17376 14116 17400 14118
rect 17456 14116 17480 14118
rect 17536 14116 17542 14118
rect 17234 14107 17542 14116
rect 17880 14074 17908 21490
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 14520 13628 14828 13637
rect 14520 13626 14526 13628
rect 14582 13626 14606 13628
rect 14662 13626 14686 13628
rect 14742 13626 14766 13628
rect 14822 13626 14828 13628
rect 14582 13574 14584 13626
rect 14764 13574 14766 13626
rect 14520 13572 14526 13574
rect 14582 13572 14606 13574
rect 14662 13572 14686 13574
rect 14742 13572 14766 13574
rect 14822 13572 14828 13574
rect 14520 13563 14828 13572
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 11806 13084 12114 13093
rect 11806 13082 11812 13084
rect 11868 13082 11892 13084
rect 11948 13082 11972 13084
rect 12028 13082 12052 13084
rect 12108 13082 12114 13084
rect 11868 13030 11870 13082
rect 12050 13030 12052 13082
rect 11806 13028 11812 13030
rect 11868 13028 11892 13030
rect 11948 13028 11972 13030
rect 12028 13028 12052 13030
rect 12108 13028 12114 13030
rect 11806 13019 12114 13028
rect 16224 12986 16252 13262
rect 16868 12986 16896 13806
rect 16948 13320 17000 13326
rect 17052 13308 17080 13874
rect 17000 13280 17080 13308
rect 16948 13262 17000 13268
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 14520 12540 14828 12549
rect 14520 12538 14526 12540
rect 14582 12538 14606 12540
rect 14662 12538 14686 12540
rect 14742 12538 14766 12540
rect 14822 12538 14828 12540
rect 14582 12486 14584 12538
rect 14764 12486 14766 12538
rect 14520 12484 14526 12486
rect 14582 12484 14606 12486
rect 14662 12484 14686 12486
rect 14742 12484 14766 12486
rect 14822 12484 14828 12486
rect 14520 12475 14828 12484
rect 16132 12442 16160 12786
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16132 12322 16160 12378
rect 16040 12294 16160 12322
rect 16040 12238 16068 12294
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16868 12170 16896 12786
rect 16960 12238 16988 13262
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17234 13084 17542 13093
rect 17234 13082 17240 13084
rect 17296 13082 17320 13084
rect 17376 13082 17400 13084
rect 17456 13082 17480 13084
rect 17536 13082 17542 13084
rect 17296 13030 17298 13082
rect 17478 13030 17480 13082
rect 17234 13028 17240 13030
rect 17296 13028 17320 13030
rect 17376 13028 17400 13030
rect 17456 13028 17480 13030
rect 17536 13028 17542 13030
rect 17234 13019 17542 13028
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 11806 11996 12114 12005
rect 11806 11994 11812 11996
rect 11868 11994 11892 11996
rect 11948 11994 11972 11996
rect 12028 11994 12052 11996
rect 12108 11994 12114 11996
rect 11868 11942 11870 11994
rect 12050 11942 12052 11994
rect 11806 11940 11812 11942
rect 11868 11940 11892 11942
rect 11948 11940 11972 11942
rect 12028 11940 12052 11942
rect 12108 11940 12114 11942
rect 11806 11931 12114 11940
rect 16868 11558 16896 12106
rect 16960 11830 16988 12174
rect 17234 11996 17542 12005
rect 17234 11994 17240 11996
rect 17296 11994 17320 11996
rect 17376 11994 17400 11996
rect 17456 11994 17480 11996
rect 17536 11994 17542 11996
rect 17296 11942 17298 11994
rect 17478 11942 17480 11994
rect 17234 11940 17240 11942
rect 17296 11940 17320 11942
rect 17376 11940 17400 11942
rect 17456 11940 17480 11942
rect 17536 11940 17542 11942
rect 17234 11931 17542 11940
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 14520 11452 14828 11461
rect 14520 11450 14526 11452
rect 14582 11450 14606 11452
rect 14662 11450 14686 11452
rect 14742 11450 14766 11452
rect 14822 11450 14828 11452
rect 14582 11398 14584 11450
rect 14764 11398 14766 11450
rect 14520 11396 14526 11398
rect 14582 11396 14606 11398
rect 14662 11396 14686 11398
rect 14742 11396 14766 11398
rect 14822 11396 14828 11398
rect 14520 11387 14828 11396
rect 16960 11354 16988 11630
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 11806 10908 12114 10917
rect 11806 10906 11812 10908
rect 11868 10906 11892 10908
rect 11948 10906 11972 10908
rect 12028 10906 12052 10908
rect 12108 10906 12114 10908
rect 11868 10854 11870 10906
rect 12050 10854 12052 10906
rect 11806 10852 11812 10854
rect 11868 10852 11892 10854
rect 11948 10852 11972 10854
rect 12028 10852 12052 10854
rect 12108 10852 12114 10854
rect 11806 10843 12114 10852
rect 17234 10908 17542 10917
rect 17234 10906 17240 10908
rect 17296 10906 17320 10908
rect 17376 10906 17400 10908
rect 17456 10906 17480 10908
rect 17536 10906 17542 10908
rect 17296 10854 17298 10906
rect 17478 10854 17480 10906
rect 17234 10852 17240 10854
rect 17296 10852 17320 10854
rect 17376 10852 17400 10854
rect 17456 10852 17480 10854
rect 17536 10852 17542 10854
rect 17234 10843 17542 10852
rect 17604 10674 17632 11698
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 14520 10364 14828 10373
rect 14520 10362 14526 10364
rect 14582 10362 14606 10364
rect 14662 10362 14686 10364
rect 14742 10362 14766 10364
rect 14822 10362 14828 10364
rect 14582 10310 14584 10362
rect 14764 10310 14766 10362
rect 14520 10308 14526 10310
rect 14582 10308 14606 10310
rect 14662 10308 14686 10310
rect 14742 10308 14766 10310
rect 14822 10308 14828 10310
rect 14520 10299 14828 10308
rect 16868 10198 16896 10406
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 16868 9926 16896 10134
rect 17236 10130 17264 10406
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17696 9926 17724 13126
rect 17880 12782 17908 14010
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 17972 12850 18000 13262
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17972 11014 18000 12786
rect 18708 12646 18736 13262
rect 19076 12850 19104 21422
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17880 10674 17908 10950
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18064 10130 18092 12038
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 6378 9820 6686 9829
rect 6378 9818 6384 9820
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6680 9818 6686 9820
rect 6440 9766 6442 9818
rect 6622 9766 6624 9818
rect 6378 9764 6384 9766
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6680 9764 6686 9766
rect 6378 9755 6686 9764
rect 11806 9820 12114 9829
rect 11806 9818 11812 9820
rect 11868 9818 11892 9820
rect 11948 9818 11972 9820
rect 12028 9818 12052 9820
rect 12108 9818 12114 9820
rect 11868 9766 11870 9818
rect 12050 9766 12052 9818
rect 11806 9764 11812 9766
rect 11868 9764 11892 9766
rect 11948 9764 11972 9766
rect 12028 9764 12052 9766
rect 12108 9764 12114 9766
rect 11806 9755 12114 9764
rect 17234 9820 17542 9829
rect 17234 9818 17240 9820
rect 17296 9818 17320 9820
rect 17376 9818 17400 9820
rect 17456 9818 17480 9820
rect 17536 9818 17542 9820
rect 17296 9766 17298 9818
rect 17478 9766 17480 9818
rect 17234 9764 17240 9766
rect 17296 9764 17320 9766
rect 17376 9764 17400 9766
rect 17456 9764 17480 9766
rect 17536 9764 17542 9766
rect 17234 9755 17542 9764
rect 18064 9722 18092 10066
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 3664 9276 3972 9285
rect 3664 9274 3670 9276
rect 3726 9274 3750 9276
rect 3806 9274 3830 9276
rect 3886 9274 3910 9276
rect 3966 9274 3972 9276
rect 3726 9222 3728 9274
rect 3908 9222 3910 9274
rect 3664 9220 3670 9222
rect 3726 9220 3750 9222
rect 3806 9220 3830 9222
rect 3886 9220 3910 9222
rect 3966 9220 3972 9222
rect 3664 9211 3972 9220
rect 9092 9276 9400 9285
rect 9092 9274 9098 9276
rect 9154 9274 9178 9276
rect 9234 9274 9258 9276
rect 9314 9274 9338 9276
rect 9394 9274 9400 9276
rect 9154 9222 9156 9274
rect 9336 9222 9338 9274
rect 9092 9220 9098 9222
rect 9154 9220 9178 9222
rect 9234 9220 9258 9222
rect 9314 9220 9338 9222
rect 9394 9220 9400 9222
rect 9092 9211 9400 9220
rect 14520 9276 14828 9285
rect 14520 9274 14526 9276
rect 14582 9274 14606 9276
rect 14662 9274 14686 9276
rect 14742 9274 14766 9276
rect 14822 9274 14828 9276
rect 14582 9222 14584 9274
rect 14764 9222 14766 9274
rect 14520 9220 14526 9222
rect 14582 9220 14606 9222
rect 14662 9220 14686 9222
rect 14742 9220 14766 9222
rect 14822 9220 14828 9222
rect 14520 9211 14828 9220
rect 6378 8732 6686 8741
rect 6378 8730 6384 8732
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6680 8730 6686 8732
rect 6440 8678 6442 8730
rect 6622 8678 6624 8730
rect 6378 8676 6384 8678
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6680 8676 6686 8678
rect 6378 8667 6686 8676
rect 11806 8732 12114 8741
rect 11806 8730 11812 8732
rect 11868 8730 11892 8732
rect 11948 8730 11972 8732
rect 12028 8730 12052 8732
rect 12108 8730 12114 8732
rect 11868 8678 11870 8730
rect 12050 8678 12052 8730
rect 11806 8676 11812 8678
rect 11868 8676 11892 8678
rect 11948 8676 11972 8678
rect 12028 8676 12052 8678
rect 12108 8676 12114 8678
rect 11806 8667 12114 8676
rect 17234 8732 17542 8741
rect 17234 8730 17240 8732
rect 17296 8730 17320 8732
rect 17376 8730 17400 8732
rect 17456 8730 17480 8732
rect 17536 8730 17542 8732
rect 17296 8678 17298 8730
rect 17478 8678 17480 8730
rect 17234 8676 17240 8678
rect 17296 8676 17320 8678
rect 17376 8676 17400 8678
rect 17456 8676 17480 8678
rect 17536 8676 17542 8678
rect 17234 8667 17542 8676
rect 3664 8188 3972 8197
rect 3664 8186 3670 8188
rect 3726 8186 3750 8188
rect 3806 8186 3830 8188
rect 3886 8186 3910 8188
rect 3966 8186 3972 8188
rect 3726 8134 3728 8186
rect 3908 8134 3910 8186
rect 3664 8132 3670 8134
rect 3726 8132 3750 8134
rect 3806 8132 3830 8134
rect 3886 8132 3910 8134
rect 3966 8132 3972 8134
rect 3664 8123 3972 8132
rect 9092 8188 9400 8197
rect 9092 8186 9098 8188
rect 9154 8186 9178 8188
rect 9234 8186 9258 8188
rect 9314 8186 9338 8188
rect 9394 8186 9400 8188
rect 9154 8134 9156 8186
rect 9336 8134 9338 8186
rect 9092 8132 9098 8134
rect 9154 8132 9178 8134
rect 9234 8132 9258 8134
rect 9314 8132 9338 8134
rect 9394 8132 9400 8134
rect 9092 8123 9400 8132
rect 14520 8188 14828 8197
rect 14520 8186 14526 8188
rect 14582 8186 14606 8188
rect 14662 8186 14686 8188
rect 14742 8186 14766 8188
rect 14822 8186 14828 8188
rect 14582 8134 14584 8186
rect 14764 8134 14766 8186
rect 14520 8132 14526 8134
rect 14582 8132 14606 8134
rect 14662 8132 14686 8134
rect 14742 8132 14766 8134
rect 14822 8132 14828 8134
rect 14520 8123 14828 8132
rect 18156 7954 18184 12582
rect 18708 12442 18736 12582
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18248 11150 18276 12378
rect 18800 12170 18828 12786
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12434 19012 12582
rect 18892 12406 19012 12434
rect 18892 12374 18920 12406
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18892 11694 18920 12310
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 9722 18644 10542
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18708 9586 18736 11086
rect 18892 10810 18920 11630
rect 18984 11626 19012 12106
rect 19076 11898 19104 12786
rect 19444 12306 19472 13126
rect 19812 12850 19840 21422
rect 19948 21244 20256 21253
rect 19948 21242 19954 21244
rect 20010 21242 20034 21244
rect 20090 21242 20114 21244
rect 20170 21242 20194 21244
rect 20250 21242 20256 21244
rect 20010 21190 20012 21242
rect 20192 21190 20194 21242
rect 19948 21188 19954 21190
rect 20010 21188 20034 21190
rect 20090 21188 20114 21190
rect 20170 21188 20194 21190
rect 20250 21188 20256 21190
rect 19948 21179 20256 21188
rect 19948 20156 20256 20165
rect 19948 20154 19954 20156
rect 20010 20154 20034 20156
rect 20090 20154 20114 20156
rect 20170 20154 20194 20156
rect 20250 20154 20256 20156
rect 20010 20102 20012 20154
rect 20192 20102 20194 20154
rect 19948 20100 19954 20102
rect 20010 20100 20034 20102
rect 20090 20100 20114 20102
rect 20170 20100 20194 20102
rect 20250 20100 20256 20102
rect 19948 20091 20256 20100
rect 19948 19068 20256 19077
rect 19948 19066 19954 19068
rect 20010 19066 20034 19068
rect 20090 19066 20114 19068
rect 20170 19066 20194 19068
rect 20250 19066 20256 19068
rect 20010 19014 20012 19066
rect 20192 19014 20194 19066
rect 19948 19012 19954 19014
rect 20010 19012 20034 19014
rect 20090 19012 20114 19014
rect 20170 19012 20194 19014
rect 20250 19012 20256 19014
rect 19948 19003 20256 19012
rect 19948 17980 20256 17989
rect 19948 17978 19954 17980
rect 20010 17978 20034 17980
rect 20090 17978 20114 17980
rect 20170 17978 20194 17980
rect 20250 17978 20256 17980
rect 20010 17926 20012 17978
rect 20192 17926 20194 17978
rect 19948 17924 19954 17926
rect 20010 17924 20034 17926
rect 20090 17924 20114 17926
rect 20170 17924 20194 17926
rect 20250 17924 20256 17926
rect 19948 17915 20256 17924
rect 19948 16892 20256 16901
rect 19948 16890 19954 16892
rect 20010 16890 20034 16892
rect 20090 16890 20114 16892
rect 20170 16890 20194 16892
rect 20250 16890 20256 16892
rect 20010 16838 20012 16890
rect 20192 16838 20194 16890
rect 19948 16836 19954 16838
rect 20010 16836 20034 16838
rect 20090 16836 20114 16838
rect 20170 16836 20194 16838
rect 20250 16836 20256 16838
rect 19948 16827 20256 16836
rect 19948 15804 20256 15813
rect 19948 15802 19954 15804
rect 20010 15802 20034 15804
rect 20090 15802 20114 15804
rect 20170 15802 20194 15804
rect 20250 15802 20256 15804
rect 20010 15750 20012 15802
rect 20192 15750 20194 15802
rect 19948 15748 19954 15750
rect 20010 15748 20034 15750
rect 20090 15748 20114 15750
rect 20170 15748 20194 15750
rect 20250 15748 20256 15750
rect 19948 15739 20256 15748
rect 19948 14716 20256 14725
rect 19948 14714 19954 14716
rect 20010 14714 20034 14716
rect 20090 14714 20114 14716
rect 20170 14714 20194 14716
rect 20250 14714 20256 14716
rect 20010 14662 20012 14714
rect 20192 14662 20194 14714
rect 19948 14660 19954 14662
rect 20010 14660 20034 14662
rect 20090 14660 20114 14662
rect 20170 14660 20194 14662
rect 20250 14660 20256 14662
rect 19948 14651 20256 14660
rect 19948 13628 20256 13637
rect 19948 13626 19954 13628
rect 20010 13626 20034 13628
rect 20090 13626 20114 13628
rect 20170 13626 20194 13628
rect 20250 13626 20256 13628
rect 20010 13574 20012 13626
rect 20192 13574 20194 13626
rect 19948 13572 19954 13574
rect 20010 13572 20034 13574
rect 20090 13572 20114 13574
rect 20170 13572 20194 13574
rect 20250 13572 20256 13574
rect 19948 13563 20256 13572
rect 20456 12850 20484 21490
rect 22662 20700 22970 20709
rect 22662 20698 22668 20700
rect 22724 20698 22748 20700
rect 22804 20698 22828 20700
rect 22884 20698 22908 20700
rect 22964 20698 22970 20700
rect 22724 20646 22726 20698
rect 22906 20646 22908 20698
rect 22662 20644 22668 20646
rect 22724 20644 22748 20646
rect 22804 20644 22828 20646
rect 22884 20644 22908 20646
rect 22964 20644 22970 20646
rect 22662 20635 22970 20644
rect 22662 19612 22970 19621
rect 22662 19610 22668 19612
rect 22724 19610 22748 19612
rect 22804 19610 22828 19612
rect 22884 19610 22908 19612
rect 22964 19610 22970 19612
rect 22724 19558 22726 19610
rect 22906 19558 22908 19610
rect 22662 19556 22668 19558
rect 22724 19556 22748 19558
rect 22804 19556 22828 19558
rect 22884 19556 22908 19558
rect 22964 19556 22970 19558
rect 22662 19547 22970 19556
rect 22662 18524 22970 18533
rect 22662 18522 22668 18524
rect 22724 18522 22748 18524
rect 22804 18522 22828 18524
rect 22884 18522 22908 18524
rect 22964 18522 22970 18524
rect 22724 18470 22726 18522
rect 22906 18470 22908 18522
rect 22662 18468 22668 18470
rect 22724 18468 22748 18470
rect 22804 18468 22828 18470
rect 22884 18468 22908 18470
rect 22964 18468 22970 18470
rect 22662 18459 22970 18468
rect 22662 17436 22970 17445
rect 22662 17434 22668 17436
rect 22724 17434 22748 17436
rect 22804 17434 22828 17436
rect 22884 17434 22908 17436
rect 22964 17434 22970 17436
rect 22724 17382 22726 17434
rect 22906 17382 22908 17434
rect 22662 17380 22668 17382
rect 22724 17380 22748 17382
rect 22804 17380 22828 17382
rect 22884 17380 22908 17382
rect 22964 17380 22970 17382
rect 22662 17371 22970 17380
rect 22662 16348 22970 16357
rect 22662 16346 22668 16348
rect 22724 16346 22748 16348
rect 22804 16346 22828 16348
rect 22884 16346 22908 16348
rect 22964 16346 22970 16348
rect 22724 16294 22726 16346
rect 22906 16294 22908 16346
rect 22662 16292 22668 16294
rect 22724 16292 22748 16294
rect 22804 16292 22828 16294
rect 22884 16292 22908 16294
rect 22964 16292 22970 16294
rect 22662 16283 22970 16292
rect 22662 15260 22970 15269
rect 22662 15258 22668 15260
rect 22724 15258 22748 15260
rect 22804 15258 22828 15260
rect 22884 15258 22908 15260
rect 22964 15258 22970 15260
rect 22724 15206 22726 15258
rect 22906 15206 22908 15258
rect 22662 15204 22668 15206
rect 22724 15204 22748 15206
rect 22804 15204 22828 15206
rect 22884 15204 22908 15206
rect 22964 15204 22970 15206
rect 22662 15195 22970 15204
rect 22662 14172 22970 14181
rect 22662 14170 22668 14172
rect 22724 14170 22748 14172
rect 22804 14170 22828 14172
rect 22884 14170 22908 14172
rect 22964 14170 22970 14172
rect 22724 14118 22726 14170
rect 22906 14118 22908 14170
rect 22662 14116 22668 14118
rect 22724 14116 22748 14118
rect 22804 14116 22828 14118
rect 22884 14116 22908 14118
rect 22964 14116 22970 14118
rect 22662 14107 22970 14116
rect 22662 13084 22970 13093
rect 22662 13082 22668 13084
rect 22724 13082 22748 13084
rect 22804 13082 22828 13084
rect 22884 13082 22908 13084
rect 22964 13082 22970 13084
rect 22724 13030 22726 13082
rect 22906 13030 22908 13082
rect 22662 13028 22668 13030
rect 22724 13028 22748 13030
rect 22804 13028 22828 13030
rect 22884 13028 22908 13030
rect 22964 13028 22970 13030
rect 22662 13019 22970 13028
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18892 10266 18920 10746
rect 18984 10674 19012 11562
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18984 10130 19012 10610
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 6378 7644 6686 7653
rect 6378 7642 6384 7644
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6680 7642 6686 7644
rect 6440 7590 6442 7642
rect 6622 7590 6624 7642
rect 6378 7588 6384 7590
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6680 7588 6686 7590
rect 6378 7579 6686 7588
rect 11806 7644 12114 7653
rect 11806 7642 11812 7644
rect 11868 7642 11892 7644
rect 11948 7642 11972 7644
rect 12028 7642 12052 7644
rect 12108 7642 12114 7644
rect 11868 7590 11870 7642
rect 12050 7590 12052 7642
rect 11806 7588 11812 7590
rect 11868 7588 11892 7590
rect 11948 7588 11972 7590
rect 12028 7588 12052 7590
rect 12108 7588 12114 7590
rect 11806 7579 12114 7588
rect 17234 7644 17542 7653
rect 17234 7642 17240 7644
rect 17296 7642 17320 7644
rect 17376 7642 17400 7644
rect 17456 7642 17480 7644
rect 17536 7642 17542 7644
rect 17296 7590 17298 7642
rect 17478 7590 17480 7642
rect 17234 7588 17240 7590
rect 17296 7588 17320 7590
rect 17376 7588 17400 7590
rect 17456 7588 17480 7590
rect 17536 7588 17542 7590
rect 17234 7579 17542 7588
rect 18064 7478 18092 7822
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18432 7342 18460 7822
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 3664 7100 3972 7109
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7035 3972 7044
rect 9092 7100 9400 7109
rect 9092 7098 9098 7100
rect 9154 7098 9178 7100
rect 9234 7098 9258 7100
rect 9314 7098 9338 7100
rect 9394 7098 9400 7100
rect 9154 7046 9156 7098
rect 9336 7046 9338 7098
rect 9092 7044 9098 7046
rect 9154 7044 9178 7046
rect 9234 7044 9258 7046
rect 9314 7044 9338 7046
rect 9394 7044 9400 7046
rect 9092 7035 9400 7044
rect 14520 7100 14828 7109
rect 14520 7098 14526 7100
rect 14582 7098 14606 7100
rect 14662 7098 14686 7100
rect 14742 7098 14766 7100
rect 14822 7098 14828 7100
rect 14582 7046 14584 7098
rect 14764 7046 14766 7098
rect 14520 7044 14526 7046
rect 14582 7044 14606 7046
rect 14662 7044 14686 7046
rect 14742 7044 14766 7046
rect 14822 7044 14828 7046
rect 14520 7035 14828 7044
rect 6378 6556 6686 6565
rect 6378 6554 6384 6556
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6680 6554 6686 6556
rect 6440 6502 6442 6554
rect 6622 6502 6624 6554
rect 6378 6500 6384 6502
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6680 6500 6686 6502
rect 6378 6491 6686 6500
rect 11806 6556 12114 6565
rect 11806 6554 11812 6556
rect 11868 6554 11892 6556
rect 11948 6554 11972 6556
rect 12028 6554 12052 6556
rect 12108 6554 12114 6556
rect 11868 6502 11870 6554
rect 12050 6502 12052 6554
rect 11806 6500 11812 6502
rect 11868 6500 11892 6502
rect 11948 6500 11972 6502
rect 12028 6500 12052 6502
rect 12108 6500 12114 6502
rect 11806 6491 12114 6500
rect 17234 6556 17542 6565
rect 17234 6554 17240 6556
rect 17296 6554 17320 6556
rect 17376 6554 17400 6556
rect 17456 6554 17480 6556
rect 17536 6554 17542 6556
rect 17296 6502 17298 6554
rect 17478 6502 17480 6554
rect 17234 6500 17240 6502
rect 17296 6500 17320 6502
rect 17376 6500 17400 6502
rect 17456 6500 17480 6502
rect 17536 6500 17542 6502
rect 17234 6491 17542 6500
rect 3664 6012 3972 6021
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5947 3972 5956
rect 9092 6012 9400 6021
rect 9092 6010 9098 6012
rect 9154 6010 9178 6012
rect 9234 6010 9258 6012
rect 9314 6010 9338 6012
rect 9394 6010 9400 6012
rect 9154 5958 9156 6010
rect 9336 5958 9338 6010
rect 9092 5956 9098 5958
rect 9154 5956 9178 5958
rect 9234 5956 9258 5958
rect 9314 5956 9338 5958
rect 9394 5956 9400 5958
rect 9092 5947 9400 5956
rect 14520 6012 14828 6021
rect 14520 6010 14526 6012
rect 14582 6010 14606 6012
rect 14662 6010 14686 6012
rect 14742 6010 14766 6012
rect 14822 6010 14828 6012
rect 14582 5958 14584 6010
rect 14764 5958 14766 6010
rect 14520 5956 14526 5958
rect 14582 5956 14606 5958
rect 14662 5956 14686 5958
rect 14742 5956 14766 5958
rect 14822 5956 14828 5958
rect 14520 5947 14828 5956
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 6378 5468 6686 5477
rect 6378 5466 6384 5468
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6680 5466 6686 5468
rect 6440 5414 6442 5466
rect 6622 5414 6624 5466
rect 6378 5412 6384 5414
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6680 5412 6686 5414
rect 6378 5403 6686 5412
rect 11806 5468 12114 5477
rect 11806 5466 11812 5468
rect 11868 5466 11892 5468
rect 11948 5466 11972 5468
rect 12028 5466 12052 5468
rect 12108 5466 12114 5468
rect 11868 5414 11870 5466
rect 12050 5414 12052 5466
rect 11806 5412 11812 5414
rect 11868 5412 11892 5414
rect 11948 5412 11972 5414
rect 12028 5412 12052 5414
rect 12108 5412 12114 5414
rect 11806 5403 12114 5412
rect 17234 5468 17542 5477
rect 17234 5466 17240 5468
rect 17296 5466 17320 5468
rect 17376 5466 17400 5468
rect 17456 5466 17480 5468
rect 17536 5466 17542 5468
rect 17296 5414 17298 5466
rect 17478 5414 17480 5466
rect 17234 5412 17240 5414
rect 17296 5412 17320 5414
rect 17376 5412 17400 5414
rect 17456 5412 17480 5414
rect 17536 5412 17542 5414
rect 17234 5403 17542 5412
rect 3664 4924 3972 4933
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4859 3972 4868
rect 9092 4924 9400 4933
rect 9092 4922 9098 4924
rect 9154 4922 9178 4924
rect 9234 4922 9258 4924
rect 9314 4922 9338 4924
rect 9394 4922 9400 4924
rect 9154 4870 9156 4922
rect 9336 4870 9338 4922
rect 9092 4868 9098 4870
rect 9154 4868 9178 4870
rect 9234 4868 9258 4870
rect 9314 4868 9338 4870
rect 9394 4868 9400 4870
rect 9092 4859 9400 4868
rect 14520 4924 14828 4933
rect 14520 4922 14526 4924
rect 14582 4922 14606 4924
rect 14662 4922 14686 4924
rect 14742 4922 14766 4924
rect 14822 4922 14828 4924
rect 14582 4870 14584 4922
rect 14764 4870 14766 4922
rect 14520 4868 14526 4870
rect 14582 4868 14606 4870
rect 14662 4868 14686 4870
rect 14742 4868 14766 4870
rect 14822 4868 14828 4870
rect 14520 4859 14828 4868
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 6378 4380 6686 4389
rect 6378 4378 6384 4380
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6680 4378 6686 4380
rect 6440 4326 6442 4378
rect 6622 4326 6624 4378
rect 6378 4324 6384 4326
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6680 4324 6686 4326
rect 6378 4315 6686 4324
rect 11806 4380 12114 4389
rect 11806 4378 11812 4380
rect 11868 4378 11892 4380
rect 11948 4378 11972 4380
rect 12028 4378 12052 4380
rect 12108 4378 12114 4380
rect 11868 4326 11870 4378
rect 12050 4326 12052 4378
rect 11806 4324 11812 4326
rect 11868 4324 11892 4326
rect 11948 4324 11972 4326
rect 12028 4324 12052 4326
rect 12108 4324 12114 4326
rect 11806 4315 12114 4324
rect 3664 3836 3972 3845
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 3664 3771 3972 3780
rect 9092 3836 9400 3845
rect 9092 3834 9098 3836
rect 9154 3834 9178 3836
rect 9234 3834 9258 3836
rect 9314 3834 9338 3836
rect 9394 3834 9400 3836
rect 9154 3782 9156 3834
rect 9336 3782 9338 3834
rect 9092 3780 9098 3782
rect 9154 3780 9178 3782
rect 9234 3780 9258 3782
rect 9314 3780 9338 3782
rect 9394 3780 9400 3782
rect 9092 3771 9400 3780
rect 14520 3836 14828 3845
rect 14520 3834 14526 3836
rect 14582 3834 14606 3836
rect 14662 3834 14686 3836
rect 14742 3834 14766 3836
rect 14822 3834 14828 3836
rect 14582 3782 14584 3834
rect 14764 3782 14766 3834
rect 14520 3780 14526 3782
rect 14582 3780 14606 3782
rect 14662 3780 14686 3782
rect 14742 3780 14766 3782
rect 14822 3780 14828 3782
rect 14520 3771 14828 3780
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 6378 3292 6686 3301
rect 6378 3290 6384 3292
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6680 3290 6686 3292
rect 6440 3238 6442 3290
rect 6622 3238 6624 3290
rect 6378 3236 6384 3238
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6680 3236 6686 3238
rect 6378 3227 6686 3236
rect 11806 3292 12114 3301
rect 11806 3290 11812 3292
rect 11868 3290 11892 3292
rect 11948 3290 11972 3292
rect 12028 3290 12052 3292
rect 12108 3290 12114 3292
rect 11868 3238 11870 3290
rect 12050 3238 12052 3290
rect 11806 3236 11812 3238
rect 11868 3236 11892 3238
rect 11948 3236 11972 3238
rect 12028 3236 12052 3238
rect 12108 3236 12114 3238
rect 11806 3227 12114 3236
rect 13004 3058 13032 3334
rect 14384 3058 14412 3334
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 3664 2748 3972 2757
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2683 3972 2692
rect 9092 2748 9400 2757
rect 9092 2746 9098 2748
rect 9154 2746 9178 2748
rect 9234 2746 9258 2748
rect 9314 2746 9338 2748
rect 9394 2746 9400 2748
rect 9154 2694 9156 2746
rect 9336 2694 9338 2746
rect 9092 2692 9098 2694
rect 9154 2692 9178 2694
rect 9234 2692 9258 2694
rect 9314 2692 9338 2694
rect 9394 2692 9400 2694
rect 9092 2683 9400 2692
rect 12360 2650 12388 2926
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 13004 2582 13032 2994
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 2056 800 2084 2382
rect 6012 800 6040 2382
rect 6378 2204 6686 2213
rect 6378 2202 6384 2204
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6680 2202 6686 2204
rect 6440 2150 6442 2202
rect 6622 2150 6624 2202
rect 6378 2148 6384 2150
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6680 2148 6686 2150
rect 6378 2139 6686 2148
rect 9968 800 9996 2382
rect 13372 2310 13400 2790
rect 14108 2650 14136 2994
rect 15672 2922 15700 4694
rect 18248 4690 18276 5510
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 17234 4380 17542 4389
rect 17234 4378 17240 4380
rect 17296 4378 17320 4380
rect 17376 4378 17400 4380
rect 17456 4378 17480 4380
rect 17536 4378 17542 4380
rect 17296 4326 17298 4378
rect 17478 4326 17480 4378
rect 17234 4324 17240 4326
rect 17296 4324 17320 4326
rect 17376 4324 17400 4326
rect 17456 4324 17480 4326
rect 17536 4324 17542 4326
rect 17234 4315 17542 4324
rect 17234 3292 17542 3301
rect 17234 3290 17240 3292
rect 17296 3290 17320 3292
rect 17376 3290 17400 3292
rect 17456 3290 17480 3292
rect 17536 3290 17542 3292
rect 17296 3238 17298 3290
rect 17478 3238 17480 3290
rect 17234 3236 17240 3238
rect 17296 3236 17320 3238
rect 17376 3236 17400 3238
rect 17456 3236 17480 3238
rect 17536 3236 17542 3238
rect 17234 3227 17542 3236
rect 18248 3126 18276 4626
rect 18432 3194 18460 7278
rect 18524 4554 18552 7686
rect 18616 4622 18644 8298
rect 18708 7818 18736 9522
rect 18892 8294 18920 9862
rect 19260 9586 19288 11018
rect 19720 10742 19748 12174
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 19720 10062 19748 10678
rect 19812 10266 19840 12786
rect 19948 12540 20256 12549
rect 19948 12538 19954 12540
rect 20010 12538 20034 12540
rect 20090 12538 20114 12540
rect 20170 12538 20194 12540
rect 20250 12538 20256 12540
rect 20010 12486 20012 12538
rect 20192 12486 20194 12538
rect 19948 12484 19954 12486
rect 20010 12484 20034 12486
rect 20090 12484 20114 12486
rect 20170 12484 20194 12486
rect 20250 12484 20256 12486
rect 19948 12475 20256 12484
rect 20456 12442 20484 12786
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 22662 11996 22970 12005
rect 22662 11994 22668 11996
rect 22724 11994 22748 11996
rect 22804 11994 22828 11996
rect 22884 11994 22908 11996
rect 22964 11994 22970 11996
rect 22724 11942 22726 11994
rect 22906 11942 22908 11994
rect 22662 11940 22668 11942
rect 22724 11940 22748 11942
rect 22804 11940 22828 11942
rect 22884 11940 22908 11942
rect 22964 11940 22970 11942
rect 22662 11931 22970 11940
rect 19948 11452 20256 11461
rect 19948 11450 19954 11452
rect 20010 11450 20034 11452
rect 20090 11450 20114 11452
rect 20170 11450 20194 11452
rect 20250 11450 20256 11452
rect 20010 11398 20012 11450
rect 20192 11398 20194 11450
rect 19948 11396 19954 11398
rect 20010 11396 20034 11398
rect 20090 11396 20114 11398
rect 20170 11396 20194 11398
rect 20250 11396 20256 11398
rect 19948 11387 20256 11396
rect 21548 11280 21600 11286
rect 21548 11222 21600 11228
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 19948 10364 20256 10373
rect 19948 10362 19954 10364
rect 20010 10362 20034 10364
rect 20090 10362 20114 10364
rect 20170 10362 20194 10364
rect 20250 10362 20256 10364
rect 20010 10310 20012 10362
rect 20192 10310 20194 10362
rect 19948 10308 19954 10310
rect 20010 10308 20034 10310
rect 20090 10308 20114 10310
rect 20170 10308 20194 10310
rect 20250 10308 20256 10310
rect 19948 10299 20256 10308
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19444 9722 19472 9998
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18892 7410 18920 7822
rect 19168 7818 19196 8434
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 19260 7546 19288 9522
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 14520 2748 14828 2757
rect 14520 2746 14526 2748
rect 14582 2746 14606 2748
rect 14662 2746 14686 2748
rect 14742 2746 14766 2748
rect 14822 2746 14828 2748
rect 14582 2694 14584 2746
rect 14764 2694 14766 2746
rect 14520 2692 14526 2694
rect 14582 2692 14606 2694
rect 14662 2692 14686 2694
rect 14742 2692 14766 2694
rect 14822 2692 14828 2694
rect 14520 2683 14828 2692
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 11806 2204 12114 2213
rect 11806 2202 11812 2204
rect 11868 2202 11892 2204
rect 11948 2202 11972 2204
rect 12028 2202 12052 2204
rect 12108 2202 12114 2204
rect 11868 2150 11870 2202
rect 12050 2150 12052 2202
rect 11806 2148 11812 2150
rect 11868 2148 11892 2150
rect 11948 2148 11972 2150
rect 12028 2148 12052 2150
rect 12108 2148 12114 2150
rect 11806 2139 12114 2148
rect 13924 800 13952 2382
rect 17234 2204 17542 2213
rect 17234 2202 17240 2204
rect 17296 2202 17320 2204
rect 17376 2202 17400 2204
rect 17456 2202 17480 2204
rect 17536 2202 17542 2204
rect 17296 2150 17298 2202
rect 17478 2150 17480 2202
rect 17234 2148 17240 2150
rect 17296 2148 17320 2150
rect 17376 2148 17400 2150
rect 17456 2148 17480 2150
rect 17536 2148 17542 2150
rect 17234 2139 17542 2148
rect 17880 800 17908 2790
rect 18892 2650 18920 7346
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5234 19380 5646
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19352 5030 19380 5170
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19352 4146 19380 4966
rect 19628 4826 19656 5578
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19536 3738 19564 4082
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19628 3534 19656 4558
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19720 2990 19748 9998
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19996 9722 20024 9930
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 21192 9586 21220 10474
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10130 21312 10406
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21376 9654 21404 10610
rect 21560 10130 21588 11222
rect 22662 10908 22970 10917
rect 22662 10906 22668 10908
rect 22724 10906 22748 10908
rect 22804 10906 22828 10908
rect 22884 10906 22908 10908
rect 22964 10906 22970 10908
rect 22724 10854 22726 10906
rect 22906 10854 22908 10906
rect 22662 10852 22668 10854
rect 22724 10852 22748 10854
rect 22804 10852 22828 10854
rect 22884 10852 22908 10854
rect 22964 10852 22970 10854
rect 22662 10843 22970 10852
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 19948 9276 20256 9285
rect 19948 9274 19954 9276
rect 20010 9274 20034 9276
rect 20090 9274 20114 9276
rect 20170 9274 20194 9276
rect 20250 9274 20256 9276
rect 20010 9222 20012 9274
rect 20192 9222 20194 9274
rect 19948 9220 19954 9222
rect 20010 9220 20034 9222
rect 20090 9220 20114 9222
rect 20170 9220 20194 9222
rect 20250 9220 20256 9222
rect 19948 9211 20256 9220
rect 20364 8498 20392 9454
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20548 8430 20576 8774
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 19948 8188 20256 8197
rect 19948 8186 19954 8188
rect 20010 8186 20034 8188
rect 20090 8186 20114 8188
rect 20170 8186 20194 8188
rect 20250 8186 20256 8188
rect 20010 8134 20012 8186
rect 20192 8134 20194 8186
rect 19948 8132 19954 8134
rect 20010 8132 20034 8134
rect 20090 8132 20114 8134
rect 20170 8132 20194 8134
rect 20250 8132 20256 8134
rect 19948 8123 20256 8132
rect 19948 7100 20256 7109
rect 19948 7098 19954 7100
rect 20010 7098 20034 7100
rect 20090 7098 20114 7100
rect 20170 7098 20194 7100
rect 20250 7098 20256 7100
rect 20010 7046 20012 7098
rect 20192 7046 20194 7098
rect 19948 7044 19954 7046
rect 20010 7044 20034 7046
rect 20090 7044 20114 7046
rect 20170 7044 20194 7046
rect 20250 7044 20256 7046
rect 19948 7035 20256 7044
rect 20456 6390 20484 8230
rect 20548 7478 20576 8366
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20444 6384 20496 6390
rect 20444 6326 20496 6332
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 19948 6012 20256 6021
rect 19948 6010 19954 6012
rect 20010 6010 20034 6012
rect 20090 6010 20114 6012
rect 20170 6010 20194 6012
rect 20250 6010 20256 6012
rect 20010 5958 20012 6010
rect 20192 5958 20194 6010
rect 19948 5956 19954 5958
rect 20010 5956 20034 5958
rect 20090 5956 20114 5958
rect 20170 5956 20194 5958
rect 20250 5956 20256 5958
rect 19948 5947 20256 5956
rect 20456 5370 20484 6054
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 19948 4924 20256 4933
rect 19948 4922 19954 4924
rect 20010 4922 20034 4924
rect 20090 4922 20114 4924
rect 20170 4922 20194 4924
rect 20250 4922 20256 4924
rect 20010 4870 20012 4922
rect 20192 4870 20194 4922
rect 19948 4868 19954 4870
rect 20010 4868 20034 4870
rect 20090 4868 20114 4870
rect 20170 4868 20194 4870
rect 20250 4868 20256 4870
rect 19948 4859 20256 4868
rect 20548 4826 20576 7414
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 19948 3836 20256 3845
rect 19948 3834 19954 3836
rect 20010 3834 20034 3836
rect 20090 3834 20114 3836
rect 20170 3834 20194 3836
rect 20250 3834 20256 3836
rect 20010 3782 20012 3834
rect 20192 3782 20194 3834
rect 19948 3780 19954 3782
rect 20010 3780 20034 3782
rect 20090 3780 20114 3782
rect 20170 3780 20194 3782
rect 20250 3780 20256 3782
rect 19948 3771 20256 3780
rect 20824 3738 20852 5238
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19948 2748 20256 2757
rect 19948 2746 19954 2748
rect 20010 2746 20034 2748
rect 20090 2746 20114 2748
rect 20170 2746 20194 2748
rect 20250 2746 20256 2748
rect 20010 2694 20012 2746
rect 20192 2694 20194 2746
rect 19948 2692 19954 2694
rect 20010 2692 20034 2694
rect 20090 2692 20114 2694
rect 20170 2692 20194 2694
rect 20250 2692 20256 2694
rect 19948 2683 20256 2692
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 20824 2446 20852 3674
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21008 2378 21036 8298
rect 21192 6458 21220 9522
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21376 3942 21404 9590
rect 21560 8294 21588 10066
rect 22662 9820 22970 9829
rect 22662 9818 22668 9820
rect 22724 9818 22748 9820
rect 22804 9818 22828 9820
rect 22884 9818 22908 9820
rect 22964 9818 22970 9820
rect 22724 9766 22726 9818
rect 22906 9766 22908 9818
rect 22662 9764 22668 9766
rect 22724 9764 22748 9766
rect 22804 9764 22828 9766
rect 22884 9764 22908 9766
rect 22964 9764 22970 9766
rect 22662 9755 22970 9764
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21652 8634 21680 8774
rect 22662 8732 22970 8741
rect 22662 8730 22668 8732
rect 22724 8730 22748 8732
rect 22804 8730 22828 8732
rect 22884 8730 22908 8732
rect 22964 8730 22970 8732
rect 22724 8678 22726 8730
rect 22906 8678 22908 8730
rect 22662 8676 22668 8678
rect 22724 8676 22748 8678
rect 22804 8676 22828 8678
rect 22884 8676 22908 8678
rect 22964 8676 22970 8678
rect 22662 8667 22970 8676
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 22662 7644 22970 7653
rect 22662 7642 22668 7644
rect 22724 7642 22748 7644
rect 22804 7642 22828 7644
rect 22884 7642 22908 7644
rect 22964 7642 22970 7644
rect 22724 7590 22726 7642
rect 22906 7590 22908 7642
rect 22662 7588 22668 7590
rect 22724 7588 22748 7590
rect 22804 7588 22828 7590
rect 22884 7588 22908 7590
rect 22964 7588 22970 7590
rect 22662 7579 22970 7588
rect 22662 6556 22970 6565
rect 22662 6554 22668 6556
rect 22724 6554 22748 6556
rect 22804 6554 22828 6556
rect 22884 6554 22908 6556
rect 22964 6554 22970 6556
rect 22724 6502 22726 6554
rect 22906 6502 22908 6554
rect 22662 6500 22668 6502
rect 22724 6500 22748 6502
rect 22804 6500 22828 6502
rect 22884 6500 22908 6502
rect 22964 6500 22970 6502
rect 22662 6491 22970 6500
rect 22662 5468 22970 5477
rect 22662 5466 22668 5468
rect 22724 5466 22748 5468
rect 22804 5466 22828 5468
rect 22884 5466 22908 5468
rect 22964 5466 22970 5468
rect 22724 5414 22726 5466
rect 22906 5414 22908 5466
rect 22662 5412 22668 5414
rect 22724 5412 22748 5414
rect 22804 5412 22828 5414
rect 22884 5412 22908 5414
rect 22964 5412 22970 5414
rect 22662 5403 22970 5412
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22008 4548 22060 4554
rect 22008 4490 22060 4496
rect 22020 4146 22048 4490
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21376 3602 21404 3878
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 20996 2372 21048 2378
rect 20996 2314 21048 2320
rect 21836 800 21864 3402
rect 22112 3194 22140 4558
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22204 3466 22232 4422
rect 22662 4380 22970 4389
rect 22662 4378 22668 4380
rect 22724 4378 22748 4380
rect 22804 4378 22828 4380
rect 22884 4378 22908 4380
rect 22964 4378 22970 4380
rect 22724 4326 22726 4378
rect 22906 4326 22908 4378
rect 22662 4324 22668 4326
rect 22724 4324 22748 4326
rect 22804 4324 22828 4326
rect 22884 4324 22908 4326
rect 22964 4324 22970 4326
rect 22662 4315 22970 4324
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22662 3292 22970 3301
rect 22662 3290 22668 3292
rect 22724 3290 22748 3292
rect 22804 3290 22828 3292
rect 22884 3290 22908 3292
rect 22964 3290 22970 3292
rect 22724 3238 22726 3290
rect 22906 3238 22908 3290
rect 22662 3236 22668 3238
rect 22724 3236 22748 3238
rect 22804 3236 22828 3238
rect 22884 3236 22908 3238
rect 22964 3236 22970 3238
rect 22662 3227 22970 3236
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 22020 2446 22048 2994
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22662 2204 22970 2213
rect 22662 2202 22668 2204
rect 22724 2202 22748 2204
rect 22804 2202 22828 2204
rect 22884 2202 22908 2204
rect 22964 2202 22970 2204
rect 22724 2150 22726 2202
rect 22906 2150 22908 2202
rect 22662 2148 22668 2150
rect 22724 2148 22748 2150
rect 22804 2148 22828 2150
rect 22884 2148 22908 2150
rect 22964 2148 22970 2150
rect 22662 2139 22970 2148
rect 2042 0 2098 800
rect 5998 0 6054 800
rect 9954 0 10010 800
rect 13910 0 13966 800
rect 17866 0 17922 800
rect 21822 0 21878 800
<< via2 >>
rect 6384 21786 6440 21788
rect 6464 21786 6520 21788
rect 6544 21786 6600 21788
rect 6624 21786 6680 21788
rect 6384 21734 6430 21786
rect 6430 21734 6440 21786
rect 6464 21734 6494 21786
rect 6494 21734 6506 21786
rect 6506 21734 6520 21786
rect 6544 21734 6558 21786
rect 6558 21734 6570 21786
rect 6570 21734 6600 21786
rect 6624 21734 6634 21786
rect 6634 21734 6680 21786
rect 6384 21732 6440 21734
rect 6464 21732 6520 21734
rect 6544 21732 6600 21734
rect 6624 21732 6680 21734
rect 11812 21786 11868 21788
rect 11892 21786 11948 21788
rect 11972 21786 12028 21788
rect 12052 21786 12108 21788
rect 11812 21734 11858 21786
rect 11858 21734 11868 21786
rect 11892 21734 11922 21786
rect 11922 21734 11934 21786
rect 11934 21734 11948 21786
rect 11972 21734 11986 21786
rect 11986 21734 11998 21786
rect 11998 21734 12028 21786
rect 12052 21734 12062 21786
rect 12062 21734 12108 21786
rect 11812 21732 11868 21734
rect 11892 21732 11948 21734
rect 11972 21732 12028 21734
rect 12052 21732 12108 21734
rect 17240 21786 17296 21788
rect 17320 21786 17376 21788
rect 17400 21786 17456 21788
rect 17480 21786 17536 21788
rect 17240 21734 17286 21786
rect 17286 21734 17296 21786
rect 17320 21734 17350 21786
rect 17350 21734 17362 21786
rect 17362 21734 17376 21786
rect 17400 21734 17414 21786
rect 17414 21734 17426 21786
rect 17426 21734 17456 21786
rect 17480 21734 17490 21786
rect 17490 21734 17536 21786
rect 17240 21732 17296 21734
rect 17320 21732 17376 21734
rect 17400 21732 17456 21734
rect 17480 21732 17536 21734
rect 22668 21786 22724 21788
rect 22748 21786 22804 21788
rect 22828 21786 22884 21788
rect 22908 21786 22964 21788
rect 22668 21734 22714 21786
rect 22714 21734 22724 21786
rect 22748 21734 22778 21786
rect 22778 21734 22790 21786
rect 22790 21734 22804 21786
rect 22828 21734 22842 21786
rect 22842 21734 22854 21786
rect 22854 21734 22884 21786
rect 22908 21734 22918 21786
rect 22918 21734 22964 21786
rect 22668 21732 22724 21734
rect 22748 21732 22804 21734
rect 22828 21732 22884 21734
rect 22908 21732 22964 21734
rect 3670 21242 3726 21244
rect 3750 21242 3806 21244
rect 3830 21242 3886 21244
rect 3910 21242 3966 21244
rect 3670 21190 3716 21242
rect 3716 21190 3726 21242
rect 3750 21190 3780 21242
rect 3780 21190 3792 21242
rect 3792 21190 3806 21242
rect 3830 21190 3844 21242
rect 3844 21190 3856 21242
rect 3856 21190 3886 21242
rect 3910 21190 3920 21242
rect 3920 21190 3966 21242
rect 3670 21188 3726 21190
rect 3750 21188 3806 21190
rect 3830 21188 3886 21190
rect 3910 21188 3966 21190
rect 3670 20154 3726 20156
rect 3750 20154 3806 20156
rect 3830 20154 3886 20156
rect 3910 20154 3966 20156
rect 3670 20102 3716 20154
rect 3716 20102 3726 20154
rect 3750 20102 3780 20154
rect 3780 20102 3792 20154
rect 3792 20102 3806 20154
rect 3830 20102 3844 20154
rect 3844 20102 3856 20154
rect 3856 20102 3886 20154
rect 3910 20102 3920 20154
rect 3920 20102 3966 20154
rect 3670 20100 3726 20102
rect 3750 20100 3806 20102
rect 3830 20100 3886 20102
rect 3910 20100 3966 20102
rect 3670 19066 3726 19068
rect 3750 19066 3806 19068
rect 3830 19066 3886 19068
rect 3910 19066 3966 19068
rect 3670 19014 3716 19066
rect 3716 19014 3726 19066
rect 3750 19014 3780 19066
rect 3780 19014 3792 19066
rect 3792 19014 3806 19066
rect 3830 19014 3844 19066
rect 3844 19014 3856 19066
rect 3856 19014 3886 19066
rect 3910 19014 3920 19066
rect 3920 19014 3966 19066
rect 3670 19012 3726 19014
rect 3750 19012 3806 19014
rect 3830 19012 3886 19014
rect 3910 19012 3966 19014
rect 3670 17978 3726 17980
rect 3750 17978 3806 17980
rect 3830 17978 3886 17980
rect 3910 17978 3966 17980
rect 3670 17926 3716 17978
rect 3716 17926 3726 17978
rect 3750 17926 3780 17978
rect 3780 17926 3792 17978
rect 3792 17926 3806 17978
rect 3830 17926 3844 17978
rect 3844 17926 3856 17978
rect 3856 17926 3886 17978
rect 3910 17926 3920 17978
rect 3920 17926 3966 17978
rect 3670 17924 3726 17926
rect 3750 17924 3806 17926
rect 3830 17924 3886 17926
rect 3910 17924 3966 17926
rect 3670 16890 3726 16892
rect 3750 16890 3806 16892
rect 3830 16890 3886 16892
rect 3910 16890 3966 16892
rect 3670 16838 3716 16890
rect 3716 16838 3726 16890
rect 3750 16838 3780 16890
rect 3780 16838 3792 16890
rect 3792 16838 3806 16890
rect 3830 16838 3844 16890
rect 3844 16838 3856 16890
rect 3856 16838 3886 16890
rect 3910 16838 3920 16890
rect 3920 16838 3966 16890
rect 3670 16836 3726 16838
rect 3750 16836 3806 16838
rect 3830 16836 3886 16838
rect 3910 16836 3966 16838
rect 3670 15802 3726 15804
rect 3750 15802 3806 15804
rect 3830 15802 3886 15804
rect 3910 15802 3966 15804
rect 3670 15750 3716 15802
rect 3716 15750 3726 15802
rect 3750 15750 3780 15802
rect 3780 15750 3792 15802
rect 3792 15750 3806 15802
rect 3830 15750 3844 15802
rect 3844 15750 3856 15802
rect 3856 15750 3886 15802
rect 3910 15750 3920 15802
rect 3920 15750 3966 15802
rect 3670 15748 3726 15750
rect 3750 15748 3806 15750
rect 3830 15748 3886 15750
rect 3910 15748 3966 15750
rect 3670 14714 3726 14716
rect 3750 14714 3806 14716
rect 3830 14714 3886 14716
rect 3910 14714 3966 14716
rect 3670 14662 3716 14714
rect 3716 14662 3726 14714
rect 3750 14662 3780 14714
rect 3780 14662 3792 14714
rect 3792 14662 3806 14714
rect 3830 14662 3844 14714
rect 3844 14662 3856 14714
rect 3856 14662 3886 14714
rect 3910 14662 3920 14714
rect 3920 14662 3966 14714
rect 3670 14660 3726 14662
rect 3750 14660 3806 14662
rect 3830 14660 3886 14662
rect 3910 14660 3966 14662
rect 3670 13626 3726 13628
rect 3750 13626 3806 13628
rect 3830 13626 3886 13628
rect 3910 13626 3966 13628
rect 3670 13574 3716 13626
rect 3716 13574 3726 13626
rect 3750 13574 3780 13626
rect 3780 13574 3792 13626
rect 3792 13574 3806 13626
rect 3830 13574 3844 13626
rect 3844 13574 3856 13626
rect 3856 13574 3886 13626
rect 3910 13574 3920 13626
rect 3920 13574 3966 13626
rect 3670 13572 3726 13574
rect 3750 13572 3806 13574
rect 3830 13572 3886 13574
rect 3910 13572 3966 13574
rect 3670 12538 3726 12540
rect 3750 12538 3806 12540
rect 3830 12538 3886 12540
rect 3910 12538 3966 12540
rect 3670 12486 3716 12538
rect 3716 12486 3726 12538
rect 3750 12486 3780 12538
rect 3780 12486 3792 12538
rect 3792 12486 3806 12538
rect 3830 12486 3844 12538
rect 3844 12486 3856 12538
rect 3856 12486 3886 12538
rect 3910 12486 3920 12538
rect 3920 12486 3966 12538
rect 3670 12484 3726 12486
rect 3750 12484 3806 12486
rect 3830 12484 3886 12486
rect 3910 12484 3966 12486
rect 6384 20698 6440 20700
rect 6464 20698 6520 20700
rect 6544 20698 6600 20700
rect 6624 20698 6680 20700
rect 6384 20646 6430 20698
rect 6430 20646 6440 20698
rect 6464 20646 6494 20698
rect 6494 20646 6506 20698
rect 6506 20646 6520 20698
rect 6544 20646 6558 20698
rect 6558 20646 6570 20698
rect 6570 20646 6600 20698
rect 6624 20646 6634 20698
rect 6634 20646 6680 20698
rect 6384 20644 6440 20646
rect 6464 20644 6520 20646
rect 6544 20644 6600 20646
rect 6624 20644 6680 20646
rect 6384 19610 6440 19612
rect 6464 19610 6520 19612
rect 6544 19610 6600 19612
rect 6624 19610 6680 19612
rect 6384 19558 6430 19610
rect 6430 19558 6440 19610
rect 6464 19558 6494 19610
rect 6494 19558 6506 19610
rect 6506 19558 6520 19610
rect 6544 19558 6558 19610
rect 6558 19558 6570 19610
rect 6570 19558 6600 19610
rect 6624 19558 6634 19610
rect 6634 19558 6680 19610
rect 6384 19556 6440 19558
rect 6464 19556 6520 19558
rect 6544 19556 6600 19558
rect 6624 19556 6680 19558
rect 6384 18522 6440 18524
rect 6464 18522 6520 18524
rect 6544 18522 6600 18524
rect 6624 18522 6680 18524
rect 6384 18470 6430 18522
rect 6430 18470 6440 18522
rect 6464 18470 6494 18522
rect 6494 18470 6506 18522
rect 6506 18470 6520 18522
rect 6544 18470 6558 18522
rect 6558 18470 6570 18522
rect 6570 18470 6600 18522
rect 6624 18470 6634 18522
rect 6634 18470 6680 18522
rect 6384 18468 6440 18470
rect 6464 18468 6520 18470
rect 6544 18468 6600 18470
rect 6624 18468 6680 18470
rect 6384 17434 6440 17436
rect 6464 17434 6520 17436
rect 6544 17434 6600 17436
rect 6624 17434 6680 17436
rect 6384 17382 6430 17434
rect 6430 17382 6440 17434
rect 6464 17382 6494 17434
rect 6494 17382 6506 17434
rect 6506 17382 6520 17434
rect 6544 17382 6558 17434
rect 6558 17382 6570 17434
rect 6570 17382 6600 17434
rect 6624 17382 6634 17434
rect 6634 17382 6680 17434
rect 6384 17380 6440 17382
rect 6464 17380 6520 17382
rect 6544 17380 6600 17382
rect 6624 17380 6680 17382
rect 6384 16346 6440 16348
rect 6464 16346 6520 16348
rect 6544 16346 6600 16348
rect 6624 16346 6680 16348
rect 6384 16294 6430 16346
rect 6430 16294 6440 16346
rect 6464 16294 6494 16346
rect 6494 16294 6506 16346
rect 6506 16294 6520 16346
rect 6544 16294 6558 16346
rect 6558 16294 6570 16346
rect 6570 16294 6600 16346
rect 6624 16294 6634 16346
rect 6634 16294 6680 16346
rect 6384 16292 6440 16294
rect 6464 16292 6520 16294
rect 6544 16292 6600 16294
rect 6624 16292 6680 16294
rect 6384 15258 6440 15260
rect 6464 15258 6520 15260
rect 6544 15258 6600 15260
rect 6624 15258 6680 15260
rect 6384 15206 6430 15258
rect 6430 15206 6440 15258
rect 6464 15206 6494 15258
rect 6494 15206 6506 15258
rect 6506 15206 6520 15258
rect 6544 15206 6558 15258
rect 6558 15206 6570 15258
rect 6570 15206 6600 15258
rect 6624 15206 6634 15258
rect 6634 15206 6680 15258
rect 6384 15204 6440 15206
rect 6464 15204 6520 15206
rect 6544 15204 6600 15206
rect 6624 15204 6680 15206
rect 6384 14170 6440 14172
rect 6464 14170 6520 14172
rect 6544 14170 6600 14172
rect 6624 14170 6680 14172
rect 6384 14118 6430 14170
rect 6430 14118 6440 14170
rect 6464 14118 6494 14170
rect 6494 14118 6506 14170
rect 6506 14118 6520 14170
rect 6544 14118 6558 14170
rect 6558 14118 6570 14170
rect 6570 14118 6600 14170
rect 6624 14118 6634 14170
rect 6634 14118 6680 14170
rect 6384 14116 6440 14118
rect 6464 14116 6520 14118
rect 6544 14116 6600 14118
rect 6624 14116 6680 14118
rect 9098 21242 9154 21244
rect 9178 21242 9234 21244
rect 9258 21242 9314 21244
rect 9338 21242 9394 21244
rect 9098 21190 9144 21242
rect 9144 21190 9154 21242
rect 9178 21190 9208 21242
rect 9208 21190 9220 21242
rect 9220 21190 9234 21242
rect 9258 21190 9272 21242
rect 9272 21190 9284 21242
rect 9284 21190 9314 21242
rect 9338 21190 9348 21242
rect 9348 21190 9394 21242
rect 9098 21188 9154 21190
rect 9178 21188 9234 21190
rect 9258 21188 9314 21190
rect 9338 21188 9394 21190
rect 9098 20154 9154 20156
rect 9178 20154 9234 20156
rect 9258 20154 9314 20156
rect 9338 20154 9394 20156
rect 9098 20102 9144 20154
rect 9144 20102 9154 20154
rect 9178 20102 9208 20154
rect 9208 20102 9220 20154
rect 9220 20102 9234 20154
rect 9258 20102 9272 20154
rect 9272 20102 9284 20154
rect 9284 20102 9314 20154
rect 9338 20102 9348 20154
rect 9348 20102 9394 20154
rect 9098 20100 9154 20102
rect 9178 20100 9234 20102
rect 9258 20100 9314 20102
rect 9338 20100 9394 20102
rect 9098 19066 9154 19068
rect 9178 19066 9234 19068
rect 9258 19066 9314 19068
rect 9338 19066 9394 19068
rect 9098 19014 9144 19066
rect 9144 19014 9154 19066
rect 9178 19014 9208 19066
rect 9208 19014 9220 19066
rect 9220 19014 9234 19066
rect 9258 19014 9272 19066
rect 9272 19014 9284 19066
rect 9284 19014 9314 19066
rect 9338 19014 9348 19066
rect 9348 19014 9394 19066
rect 9098 19012 9154 19014
rect 9178 19012 9234 19014
rect 9258 19012 9314 19014
rect 9338 19012 9394 19014
rect 9098 17978 9154 17980
rect 9178 17978 9234 17980
rect 9258 17978 9314 17980
rect 9338 17978 9394 17980
rect 9098 17926 9144 17978
rect 9144 17926 9154 17978
rect 9178 17926 9208 17978
rect 9208 17926 9220 17978
rect 9220 17926 9234 17978
rect 9258 17926 9272 17978
rect 9272 17926 9284 17978
rect 9284 17926 9314 17978
rect 9338 17926 9348 17978
rect 9348 17926 9394 17978
rect 9098 17924 9154 17926
rect 9178 17924 9234 17926
rect 9258 17924 9314 17926
rect 9338 17924 9394 17926
rect 9098 16890 9154 16892
rect 9178 16890 9234 16892
rect 9258 16890 9314 16892
rect 9338 16890 9394 16892
rect 9098 16838 9144 16890
rect 9144 16838 9154 16890
rect 9178 16838 9208 16890
rect 9208 16838 9220 16890
rect 9220 16838 9234 16890
rect 9258 16838 9272 16890
rect 9272 16838 9284 16890
rect 9284 16838 9314 16890
rect 9338 16838 9348 16890
rect 9348 16838 9394 16890
rect 9098 16836 9154 16838
rect 9178 16836 9234 16838
rect 9258 16836 9314 16838
rect 9338 16836 9394 16838
rect 9098 15802 9154 15804
rect 9178 15802 9234 15804
rect 9258 15802 9314 15804
rect 9338 15802 9394 15804
rect 9098 15750 9144 15802
rect 9144 15750 9154 15802
rect 9178 15750 9208 15802
rect 9208 15750 9220 15802
rect 9220 15750 9234 15802
rect 9258 15750 9272 15802
rect 9272 15750 9284 15802
rect 9284 15750 9314 15802
rect 9338 15750 9348 15802
rect 9348 15750 9394 15802
rect 9098 15748 9154 15750
rect 9178 15748 9234 15750
rect 9258 15748 9314 15750
rect 9338 15748 9394 15750
rect 9098 14714 9154 14716
rect 9178 14714 9234 14716
rect 9258 14714 9314 14716
rect 9338 14714 9394 14716
rect 9098 14662 9144 14714
rect 9144 14662 9154 14714
rect 9178 14662 9208 14714
rect 9208 14662 9220 14714
rect 9220 14662 9234 14714
rect 9258 14662 9272 14714
rect 9272 14662 9284 14714
rect 9284 14662 9314 14714
rect 9338 14662 9348 14714
rect 9348 14662 9394 14714
rect 9098 14660 9154 14662
rect 9178 14660 9234 14662
rect 9258 14660 9314 14662
rect 9338 14660 9394 14662
rect 9098 13626 9154 13628
rect 9178 13626 9234 13628
rect 9258 13626 9314 13628
rect 9338 13626 9394 13628
rect 9098 13574 9144 13626
rect 9144 13574 9154 13626
rect 9178 13574 9208 13626
rect 9208 13574 9220 13626
rect 9220 13574 9234 13626
rect 9258 13574 9272 13626
rect 9272 13574 9284 13626
rect 9284 13574 9314 13626
rect 9338 13574 9348 13626
rect 9348 13574 9394 13626
rect 9098 13572 9154 13574
rect 9178 13572 9234 13574
rect 9258 13572 9314 13574
rect 9338 13572 9394 13574
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6430 13082
rect 6430 13030 6440 13082
rect 6464 13030 6494 13082
rect 6494 13030 6506 13082
rect 6506 13030 6520 13082
rect 6544 13030 6558 13082
rect 6558 13030 6570 13082
rect 6570 13030 6600 13082
rect 6624 13030 6634 13082
rect 6634 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 9098 12538 9154 12540
rect 9178 12538 9234 12540
rect 9258 12538 9314 12540
rect 9338 12538 9394 12540
rect 9098 12486 9144 12538
rect 9144 12486 9154 12538
rect 9178 12486 9208 12538
rect 9208 12486 9220 12538
rect 9220 12486 9234 12538
rect 9258 12486 9272 12538
rect 9272 12486 9284 12538
rect 9284 12486 9314 12538
rect 9338 12486 9348 12538
rect 9348 12486 9394 12538
rect 9098 12484 9154 12486
rect 9178 12484 9234 12486
rect 9258 12484 9314 12486
rect 9338 12484 9394 12486
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6430 11994
rect 6430 11942 6440 11994
rect 6464 11942 6494 11994
rect 6494 11942 6506 11994
rect 6506 11942 6520 11994
rect 6544 11942 6558 11994
rect 6558 11942 6570 11994
rect 6570 11942 6600 11994
rect 6624 11942 6634 11994
rect 6634 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 3670 11450 3726 11452
rect 3750 11450 3806 11452
rect 3830 11450 3886 11452
rect 3910 11450 3966 11452
rect 3670 11398 3716 11450
rect 3716 11398 3726 11450
rect 3750 11398 3780 11450
rect 3780 11398 3792 11450
rect 3792 11398 3806 11450
rect 3830 11398 3844 11450
rect 3844 11398 3856 11450
rect 3856 11398 3886 11450
rect 3910 11398 3920 11450
rect 3920 11398 3966 11450
rect 3670 11396 3726 11398
rect 3750 11396 3806 11398
rect 3830 11396 3886 11398
rect 3910 11396 3966 11398
rect 9098 11450 9154 11452
rect 9178 11450 9234 11452
rect 9258 11450 9314 11452
rect 9338 11450 9394 11452
rect 9098 11398 9144 11450
rect 9144 11398 9154 11450
rect 9178 11398 9208 11450
rect 9208 11398 9220 11450
rect 9220 11398 9234 11450
rect 9258 11398 9272 11450
rect 9272 11398 9284 11450
rect 9284 11398 9314 11450
rect 9338 11398 9348 11450
rect 9348 11398 9394 11450
rect 9098 11396 9154 11398
rect 9178 11396 9234 11398
rect 9258 11396 9314 11398
rect 9338 11396 9394 11398
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6430 10906
rect 6430 10854 6440 10906
rect 6464 10854 6494 10906
rect 6494 10854 6506 10906
rect 6506 10854 6520 10906
rect 6544 10854 6558 10906
rect 6558 10854 6570 10906
rect 6570 10854 6600 10906
rect 6624 10854 6634 10906
rect 6634 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 3670 10362 3726 10364
rect 3750 10362 3806 10364
rect 3830 10362 3886 10364
rect 3910 10362 3966 10364
rect 3670 10310 3716 10362
rect 3716 10310 3726 10362
rect 3750 10310 3780 10362
rect 3780 10310 3792 10362
rect 3792 10310 3806 10362
rect 3830 10310 3844 10362
rect 3844 10310 3856 10362
rect 3856 10310 3886 10362
rect 3910 10310 3920 10362
rect 3920 10310 3966 10362
rect 3670 10308 3726 10310
rect 3750 10308 3806 10310
rect 3830 10308 3886 10310
rect 3910 10308 3966 10310
rect 9098 10362 9154 10364
rect 9178 10362 9234 10364
rect 9258 10362 9314 10364
rect 9338 10362 9394 10364
rect 9098 10310 9144 10362
rect 9144 10310 9154 10362
rect 9178 10310 9208 10362
rect 9208 10310 9220 10362
rect 9220 10310 9234 10362
rect 9258 10310 9272 10362
rect 9272 10310 9284 10362
rect 9284 10310 9314 10362
rect 9338 10310 9348 10362
rect 9348 10310 9394 10362
rect 9098 10308 9154 10310
rect 9178 10308 9234 10310
rect 9258 10308 9314 10310
rect 9338 10308 9394 10310
rect 14526 21242 14582 21244
rect 14606 21242 14662 21244
rect 14686 21242 14742 21244
rect 14766 21242 14822 21244
rect 14526 21190 14572 21242
rect 14572 21190 14582 21242
rect 14606 21190 14636 21242
rect 14636 21190 14648 21242
rect 14648 21190 14662 21242
rect 14686 21190 14700 21242
rect 14700 21190 14712 21242
rect 14712 21190 14742 21242
rect 14766 21190 14776 21242
rect 14776 21190 14822 21242
rect 14526 21188 14582 21190
rect 14606 21188 14662 21190
rect 14686 21188 14742 21190
rect 14766 21188 14822 21190
rect 11812 20698 11868 20700
rect 11892 20698 11948 20700
rect 11972 20698 12028 20700
rect 12052 20698 12108 20700
rect 11812 20646 11858 20698
rect 11858 20646 11868 20698
rect 11892 20646 11922 20698
rect 11922 20646 11934 20698
rect 11934 20646 11948 20698
rect 11972 20646 11986 20698
rect 11986 20646 11998 20698
rect 11998 20646 12028 20698
rect 12052 20646 12062 20698
rect 12062 20646 12108 20698
rect 11812 20644 11868 20646
rect 11892 20644 11948 20646
rect 11972 20644 12028 20646
rect 12052 20644 12108 20646
rect 17240 20698 17296 20700
rect 17320 20698 17376 20700
rect 17400 20698 17456 20700
rect 17480 20698 17536 20700
rect 17240 20646 17286 20698
rect 17286 20646 17296 20698
rect 17320 20646 17350 20698
rect 17350 20646 17362 20698
rect 17362 20646 17376 20698
rect 17400 20646 17414 20698
rect 17414 20646 17426 20698
rect 17426 20646 17456 20698
rect 17480 20646 17490 20698
rect 17490 20646 17536 20698
rect 17240 20644 17296 20646
rect 17320 20644 17376 20646
rect 17400 20644 17456 20646
rect 17480 20644 17536 20646
rect 14526 20154 14582 20156
rect 14606 20154 14662 20156
rect 14686 20154 14742 20156
rect 14766 20154 14822 20156
rect 14526 20102 14572 20154
rect 14572 20102 14582 20154
rect 14606 20102 14636 20154
rect 14636 20102 14648 20154
rect 14648 20102 14662 20154
rect 14686 20102 14700 20154
rect 14700 20102 14712 20154
rect 14712 20102 14742 20154
rect 14766 20102 14776 20154
rect 14776 20102 14822 20154
rect 14526 20100 14582 20102
rect 14606 20100 14662 20102
rect 14686 20100 14742 20102
rect 14766 20100 14822 20102
rect 11812 19610 11868 19612
rect 11892 19610 11948 19612
rect 11972 19610 12028 19612
rect 12052 19610 12108 19612
rect 11812 19558 11858 19610
rect 11858 19558 11868 19610
rect 11892 19558 11922 19610
rect 11922 19558 11934 19610
rect 11934 19558 11948 19610
rect 11972 19558 11986 19610
rect 11986 19558 11998 19610
rect 11998 19558 12028 19610
rect 12052 19558 12062 19610
rect 12062 19558 12108 19610
rect 11812 19556 11868 19558
rect 11892 19556 11948 19558
rect 11972 19556 12028 19558
rect 12052 19556 12108 19558
rect 17240 19610 17296 19612
rect 17320 19610 17376 19612
rect 17400 19610 17456 19612
rect 17480 19610 17536 19612
rect 17240 19558 17286 19610
rect 17286 19558 17296 19610
rect 17320 19558 17350 19610
rect 17350 19558 17362 19610
rect 17362 19558 17376 19610
rect 17400 19558 17414 19610
rect 17414 19558 17426 19610
rect 17426 19558 17456 19610
rect 17480 19558 17490 19610
rect 17490 19558 17536 19610
rect 17240 19556 17296 19558
rect 17320 19556 17376 19558
rect 17400 19556 17456 19558
rect 17480 19556 17536 19558
rect 14526 19066 14582 19068
rect 14606 19066 14662 19068
rect 14686 19066 14742 19068
rect 14766 19066 14822 19068
rect 14526 19014 14572 19066
rect 14572 19014 14582 19066
rect 14606 19014 14636 19066
rect 14636 19014 14648 19066
rect 14648 19014 14662 19066
rect 14686 19014 14700 19066
rect 14700 19014 14712 19066
rect 14712 19014 14742 19066
rect 14766 19014 14776 19066
rect 14776 19014 14822 19066
rect 14526 19012 14582 19014
rect 14606 19012 14662 19014
rect 14686 19012 14742 19014
rect 14766 19012 14822 19014
rect 11812 18522 11868 18524
rect 11892 18522 11948 18524
rect 11972 18522 12028 18524
rect 12052 18522 12108 18524
rect 11812 18470 11858 18522
rect 11858 18470 11868 18522
rect 11892 18470 11922 18522
rect 11922 18470 11934 18522
rect 11934 18470 11948 18522
rect 11972 18470 11986 18522
rect 11986 18470 11998 18522
rect 11998 18470 12028 18522
rect 12052 18470 12062 18522
rect 12062 18470 12108 18522
rect 11812 18468 11868 18470
rect 11892 18468 11948 18470
rect 11972 18468 12028 18470
rect 12052 18468 12108 18470
rect 17240 18522 17296 18524
rect 17320 18522 17376 18524
rect 17400 18522 17456 18524
rect 17480 18522 17536 18524
rect 17240 18470 17286 18522
rect 17286 18470 17296 18522
rect 17320 18470 17350 18522
rect 17350 18470 17362 18522
rect 17362 18470 17376 18522
rect 17400 18470 17414 18522
rect 17414 18470 17426 18522
rect 17426 18470 17456 18522
rect 17480 18470 17490 18522
rect 17490 18470 17536 18522
rect 17240 18468 17296 18470
rect 17320 18468 17376 18470
rect 17400 18468 17456 18470
rect 17480 18468 17536 18470
rect 14526 17978 14582 17980
rect 14606 17978 14662 17980
rect 14686 17978 14742 17980
rect 14766 17978 14822 17980
rect 14526 17926 14572 17978
rect 14572 17926 14582 17978
rect 14606 17926 14636 17978
rect 14636 17926 14648 17978
rect 14648 17926 14662 17978
rect 14686 17926 14700 17978
rect 14700 17926 14712 17978
rect 14712 17926 14742 17978
rect 14766 17926 14776 17978
rect 14776 17926 14822 17978
rect 14526 17924 14582 17926
rect 14606 17924 14662 17926
rect 14686 17924 14742 17926
rect 14766 17924 14822 17926
rect 11812 17434 11868 17436
rect 11892 17434 11948 17436
rect 11972 17434 12028 17436
rect 12052 17434 12108 17436
rect 11812 17382 11858 17434
rect 11858 17382 11868 17434
rect 11892 17382 11922 17434
rect 11922 17382 11934 17434
rect 11934 17382 11948 17434
rect 11972 17382 11986 17434
rect 11986 17382 11998 17434
rect 11998 17382 12028 17434
rect 12052 17382 12062 17434
rect 12062 17382 12108 17434
rect 11812 17380 11868 17382
rect 11892 17380 11948 17382
rect 11972 17380 12028 17382
rect 12052 17380 12108 17382
rect 17240 17434 17296 17436
rect 17320 17434 17376 17436
rect 17400 17434 17456 17436
rect 17480 17434 17536 17436
rect 17240 17382 17286 17434
rect 17286 17382 17296 17434
rect 17320 17382 17350 17434
rect 17350 17382 17362 17434
rect 17362 17382 17376 17434
rect 17400 17382 17414 17434
rect 17414 17382 17426 17434
rect 17426 17382 17456 17434
rect 17480 17382 17490 17434
rect 17490 17382 17536 17434
rect 17240 17380 17296 17382
rect 17320 17380 17376 17382
rect 17400 17380 17456 17382
rect 17480 17380 17536 17382
rect 14526 16890 14582 16892
rect 14606 16890 14662 16892
rect 14686 16890 14742 16892
rect 14766 16890 14822 16892
rect 14526 16838 14572 16890
rect 14572 16838 14582 16890
rect 14606 16838 14636 16890
rect 14636 16838 14648 16890
rect 14648 16838 14662 16890
rect 14686 16838 14700 16890
rect 14700 16838 14712 16890
rect 14712 16838 14742 16890
rect 14766 16838 14776 16890
rect 14776 16838 14822 16890
rect 14526 16836 14582 16838
rect 14606 16836 14662 16838
rect 14686 16836 14742 16838
rect 14766 16836 14822 16838
rect 11812 16346 11868 16348
rect 11892 16346 11948 16348
rect 11972 16346 12028 16348
rect 12052 16346 12108 16348
rect 11812 16294 11858 16346
rect 11858 16294 11868 16346
rect 11892 16294 11922 16346
rect 11922 16294 11934 16346
rect 11934 16294 11948 16346
rect 11972 16294 11986 16346
rect 11986 16294 11998 16346
rect 11998 16294 12028 16346
rect 12052 16294 12062 16346
rect 12062 16294 12108 16346
rect 11812 16292 11868 16294
rect 11892 16292 11948 16294
rect 11972 16292 12028 16294
rect 12052 16292 12108 16294
rect 17240 16346 17296 16348
rect 17320 16346 17376 16348
rect 17400 16346 17456 16348
rect 17480 16346 17536 16348
rect 17240 16294 17286 16346
rect 17286 16294 17296 16346
rect 17320 16294 17350 16346
rect 17350 16294 17362 16346
rect 17362 16294 17376 16346
rect 17400 16294 17414 16346
rect 17414 16294 17426 16346
rect 17426 16294 17456 16346
rect 17480 16294 17490 16346
rect 17490 16294 17536 16346
rect 17240 16292 17296 16294
rect 17320 16292 17376 16294
rect 17400 16292 17456 16294
rect 17480 16292 17536 16294
rect 14526 15802 14582 15804
rect 14606 15802 14662 15804
rect 14686 15802 14742 15804
rect 14766 15802 14822 15804
rect 14526 15750 14572 15802
rect 14572 15750 14582 15802
rect 14606 15750 14636 15802
rect 14636 15750 14648 15802
rect 14648 15750 14662 15802
rect 14686 15750 14700 15802
rect 14700 15750 14712 15802
rect 14712 15750 14742 15802
rect 14766 15750 14776 15802
rect 14776 15750 14822 15802
rect 14526 15748 14582 15750
rect 14606 15748 14662 15750
rect 14686 15748 14742 15750
rect 14766 15748 14822 15750
rect 11812 15258 11868 15260
rect 11892 15258 11948 15260
rect 11972 15258 12028 15260
rect 12052 15258 12108 15260
rect 11812 15206 11858 15258
rect 11858 15206 11868 15258
rect 11892 15206 11922 15258
rect 11922 15206 11934 15258
rect 11934 15206 11948 15258
rect 11972 15206 11986 15258
rect 11986 15206 11998 15258
rect 11998 15206 12028 15258
rect 12052 15206 12062 15258
rect 12062 15206 12108 15258
rect 11812 15204 11868 15206
rect 11892 15204 11948 15206
rect 11972 15204 12028 15206
rect 12052 15204 12108 15206
rect 17240 15258 17296 15260
rect 17320 15258 17376 15260
rect 17400 15258 17456 15260
rect 17480 15258 17536 15260
rect 17240 15206 17286 15258
rect 17286 15206 17296 15258
rect 17320 15206 17350 15258
rect 17350 15206 17362 15258
rect 17362 15206 17376 15258
rect 17400 15206 17414 15258
rect 17414 15206 17426 15258
rect 17426 15206 17456 15258
rect 17480 15206 17490 15258
rect 17490 15206 17536 15258
rect 17240 15204 17296 15206
rect 17320 15204 17376 15206
rect 17400 15204 17456 15206
rect 17480 15204 17536 15206
rect 14526 14714 14582 14716
rect 14606 14714 14662 14716
rect 14686 14714 14742 14716
rect 14766 14714 14822 14716
rect 14526 14662 14572 14714
rect 14572 14662 14582 14714
rect 14606 14662 14636 14714
rect 14636 14662 14648 14714
rect 14648 14662 14662 14714
rect 14686 14662 14700 14714
rect 14700 14662 14712 14714
rect 14712 14662 14742 14714
rect 14766 14662 14776 14714
rect 14776 14662 14822 14714
rect 14526 14660 14582 14662
rect 14606 14660 14662 14662
rect 14686 14660 14742 14662
rect 14766 14660 14822 14662
rect 11812 14170 11868 14172
rect 11892 14170 11948 14172
rect 11972 14170 12028 14172
rect 12052 14170 12108 14172
rect 11812 14118 11858 14170
rect 11858 14118 11868 14170
rect 11892 14118 11922 14170
rect 11922 14118 11934 14170
rect 11934 14118 11948 14170
rect 11972 14118 11986 14170
rect 11986 14118 11998 14170
rect 11998 14118 12028 14170
rect 12052 14118 12062 14170
rect 12062 14118 12108 14170
rect 11812 14116 11868 14118
rect 11892 14116 11948 14118
rect 11972 14116 12028 14118
rect 12052 14116 12108 14118
rect 17240 14170 17296 14172
rect 17320 14170 17376 14172
rect 17400 14170 17456 14172
rect 17480 14170 17536 14172
rect 17240 14118 17286 14170
rect 17286 14118 17296 14170
rect 17320 14118 17350 14170
rect 17350 14118 17362 14170
rect 17362 14118 17376 14170
rect 17400 14118 17414 14170
rect 17414 14118 17426 14170
rect 17426 14118 17456 14170
rect 17480 14118 17490 14170
rect 17490 14118 17536 14170
rect 17240 14116 17296 14118
rect 17320 14116 17376 14118
rect 17400 14116 17456 14118
rect 17480 14116 17536 14118
rect 14526 13626 14582 13628
rect 14606 13626 14662 13628
rect 14686 13626 14742 13628
rect 14766 13626 14822 13628
rect 14526 13574 14572 13626
rect 14572 13574 14582 13626
rect 14606 13574 14636 13626
rect 14636 13574 14648 13626
rect 14648 13574 14662 13626
rect 14686 13574 14700 13626
rect 14700 13574 14712 13626
rect 14712 13574 14742 13626
rect 14766 13574 14776 13626
rect 14776 13574 14822 13626
rect 14526 13572 14582 13574
rect 14606 13572 14662 13574
rect 14686 13572 14742 13574
rect 14766 13572 14822 13574
rect 11812 13082 11868 13084
rect 11892 13082 11948 13084
rect 11972 13082 12028 13084
rect 12052 13082 12108 13084
rect 11812 13030 11858 13082
rect 11858 13030 11868 13082
rect 11892 13030 11922 13082
rect 11922 13030 11934 13082
rect 11934 13030 11948 13082
rect 11972 13030 11986 13082
rect 11986 13030 11998 13082
rect 11998 13030 12028 13082
rect 12052 13030 12062 13082
rect 12062 13030 12108 13082
rect 11812 13028 11868 13030
rect 11892 13028 11948 13030
rect 11972 13028 12028 13030
rect 12052 13028 12108 13030
rect 14526 12538 14582 12540
rect 14606 12538 14662 12540
rect 14686 12538 14742 12540
rect 14766 12538 14822 12540
rect 14526 12486 14572 12538
rect 14572 12486 14582 12538
rect 14606 12486 14636 12538
rect 14636 12486 14648 12538
rect 14648 12486 14662 12538
rect 14686 12486 14700 12538
rect 14700 12486 14712 12538
rect 14712 12486 14742 12538
rect 14766 12486 14776 12538
rect 14776 12486 14822 12538
rect 14526 12484 14582 12486
rect 14606 12484 14662 12486
rect 14686 12484 14742 12486
rect 14766 12484 14822 12486
rect 17240 13082 17296 13084
rect 17320 13082 17376 13084
rect 17400 13082 17456 13084
rect 17480 13082 17536 13084
rect 17240 13030 17286 13082
rect 17286 13030 17296 13082
rect 17320 13030 17350 13082
rect 17350 13030 17362 13082
rect 17362 13030 17376 13082
rect 17400 13030 17414 13082
rect 17414 13030 17426 13082
rect 17426 13030 17456 13082
rect 17480 13030 17490 13082
rect 17490 13030 17536 13082
rect 17240 13028 17296 13030
rect 17320 13028 17376 13030
rect 17400 13028 17456 13030
rect 17480 13028 17536 13030
rect 11812 11994 11868 11996
rect 11892 11994 11948 11996
rect 11972 11994 12028 11996
rect 12052 11994 12108 11996
rect 11812 11942 11858 11994
rect 11858 11942 11868 11994
rect 11892 11942 11922 11994
rect 11922 11942 11934 11994
rect 11934 11942 11948 11994
rect 11972 11942 11986 11994
rect 11986 11942 11998 11994
rect 11998 11942 12028 11994
rect 12052 11942 12062 11994
rect 12062 11942 12108 11994
rect 11812 11940 11868 11942
rect 11892 11940 11948 11942
rect 11972 11940 12028 11942
rect 12052 11940 12108 11942
rect 17240 11994 17296 11996
rect 17320 11994 17376 11996
rect 17400 11994 17456 11996
rect 17480 11994 17536 11996
rect 17240 11942 17286 11994
rect 17286 11942 17296 11994
rect 17320 11942 17350 11994
rect 17350 11942 17362 11994
rect 17362 11942 17376 11994
rect 17400 11942 17414 11994
rect 17414 11942 17426 11994
rect 17426 11942 17456 11994
rect 17480 11942 17490 11994
rect 17490 11942 17536 11994
rect 17240 11940 17296 11942
rect 17320 11940 17376 11942
rect 17400 11940 17456 11942
rect 17480 11940 17536 11942
rect 14526 11450 14582 11452
rect 14606 11450 14662 11452
rect 14686 11450 14742 11452
rect 14766 11450 14822 11452
rect 14526 11398 14572 11450
rect 14572 11398 14582 11450
rect 14606 11398 14636 11450
rect 14636 11398 14648 11450
rect 14648 11398 14662 11450
rect 14686 11398 14700 11450
rect 14700 11398 14712 11450
rect 14712 11398 14742 11450
rect 14766 11398 14776 11450
rect 14776 11398 14822 11450
rect 14526 11396 14582 11398
rect 14606 11396 14662 11398
rect 14686 11396 14742 11398
rect 14766 11396 14822 11398
rect 11812 10906 11868 10908
rect 11892 10906 11948 10908
rect 11972 10906 12028 10908
rect 12052 10906 12108 10908
rect 11812 10854 11858 10906
rect 11858 10854 11868 10906
rect 11892 10854 11922 10906
rect 11922 10854 11934 10906
rect 11934 10854 11948 10906
rect 11972 10854 11986 10906
rect 11986 10854 11998 10906
rect 11998 10854 12028 10906
rect 12052 10854 12062 10906
rect 12062 10854 12108 10906
rect 11812 10852 11868 10854
rect 11892 10852 11948 10854
rect 11972 10852 12028 10854
rect 12052 10852 12108 10854
rect 17240 10906 17296 10908
rect 17320 10906 17376 10908
rect 17400 10906 17456 10908
rect 17480 10906 17536 10908
rect 17240 10854 17286 10906
rect 17286 10854 17296 10906
rect 17320 10854 17350 10906
rect 17350 10854 17362 10906
rect 17362 10854 17376 10906
rect 17400 10854 17414 10906
rect 17414 10854 17426 10906
rect 17426 10854 17456 10906
rect 17480 10854 17490 10906
rect 17490 10854 17536 10906
rect 17240 10852 17296 10854
rect 17320 10852 17376 10854
rect 17400 10852 17456 10854
rect 17480 10852 17536 10854
rect 14526 10362 14582 10364
rect 14606 10362 14662 10364
rect 14686 10362 14742 10364
rect 14766 10362 14822 10364
rect 14526 10310 14572 10362
rect 14572 10310 14582 10362
rect 14606 10310 14636 10362
rect 14636 10310 14648 10362
rect 14648 10310 14662 10362
rect 14686 10310 14700 10362
rect 14700 10310 14712 10362
rect 14712 10310 14742 10362
rect 14766 10310 14776 10362
rect 14776 10310 14822 10362
rect 14526 10308 14582 10310
rect 14606 10308 14662 10310
rect 14686 10308 14742 10310
rect 14766 10308 14822 10310
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6430 9818
rect 6430 9766 6440 9818
rect 6464 9766 6494 9818
rect 6494 9766 6506 9818
rect 6506 9766 6520 9818
rect 6544 9766 6558 9818
rect 6558 9766 6570 9818
rect 6570 9766 6600 9818
rect 6624 9766 6634 9818
rect 6634 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 11812 9818 11868 9820
rect 11892 9818 11948 9820
rect 11972 9818 12028 9820
rect 12052 9818 12108 9820
rect 11812 9766 11858 9818
rect 11858 9766 11868 9818
rect 11892 9766 11922 9818
rect 11922 9766 11934 9818
rect 11934 9766 11948 9818
rect 11972 9766 11986 9818
rect 11986 9766 11998 9818
rect 11998 9766 12028 9818
rect 12052 9766 12062 9818
rect 12062 9766 12108 9818
rect 11812 9764 11868 9766
rect 11892 9764 11948 9766
rect 11972 9764 12028 9766
rect 12052 9764 12108 9766
rect 17240 9818 17296 9820
rect 17320 9818 17376 9820
rect 17400 9818 17456 9820
rect 17480 9818 17536 9820
rect 17240 9766 17286 9818
rect 17286 9766 17296 9818
rect 17320 9766 17350 9818
rect 17350 9766 17362 9818
rect 17362 9766 17376 9818
rect 17400 9766 17414 9818
rect 17414 9766 17426 9818
rect 17426 9766 17456 9818
rect 17480 9766 17490 9818
rect 17490 9766 17536 9818
rect 17240 9764 17296 9766
rect 17320 9764 17376 9766
rect 17400 9764 17456 9766
rect 17480 9764 17536 9766
rect 3670 9274 3726 9276
rect 3750 9274 3806 9276
rect 3830 9274 3886 9276
rect 3910 9274 3966 9276
rect 3670 9222 3716 9274
rect 3716 9222 3726 9274
rect 3750 9222 3780 9274
rect 3780 9222 3792 9274
rect 3792 9222 3806 9274
rect 3830 9222 3844 9274
rect 3844 9222 3856 9274
rect 3856 9222 3886 9274
rect 3910 9222 3920 9274
rect 3920 9222 3966 9274
rect 3670 9220 3726 9222
rect 3750 9220 3806 9222
rect 3830 9220 3886 9222
rect 3910 9220 3966 9222
rect 9098 9274 9154 9276
rect 9178 9274 9234 9276
rect 9258 9274 9314 9276
rect 9338 9274 9394 9276
rect 9098 9222 9144 9274
rect 9144 9222 9154 9274
rect 9178 9222 9208 9274
rect 9208 9222 9220 9274
rect 9220 9222 9234 9274
rect 9258 9222 9272 9274
rect 9272 9222 9284 9274
rect 9284 9222 9314 9274
rect 9338 9222 9348 9274
rect 9348 9222 9394 9274
rect 9098 9220 9154 9222
rect 9178 9220 9234 9222
rect 9258 9220 9314 9222
rect 9338 9220 9394 9222
rect 14526 9274 14582 9276
rect 14606 9274 14662 9276
rect 14686 9274 14742 9276
rect 14766 9274 14822 9276
rect 14526 9222 14572 9274
rect 14572 9222 14582 9274
rect 14606 9222 14636 9274
rect 14636 9222 14648 9274
rect 14648 9222 14662 9274
rect 14686 9222 14700 9274
rect 14700 9222 14712 9274
rect 14712 9222 14742 9274
rect 14766 9222 14776 9274
rect 14776 9222 14822 9274
rect 14526 9220 14582 9222
rect 14606 9220 14662 9222
rect 14686 9220 14742 9222
rect 14766 9220 14822 9222
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6430 8730
rect 6430 8678 6440 8730
rect 6464 8678 6494 8730
rect 6494 8678 6506 8730
rect 6506 8678 6520 8730
rect 6544 8678 6558 8730
rect 6558 8678 6570 8730
rect 6570 8678 6600 8730
rect 6624 8678 6634 8730
rect 6634 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 11812 8730 11868 8732
rect 11892 8730 11948 8732
rect 11972 8730 12028 8732
rect 12052 8730 12108 8732
rect 11812 8678 11858 8730
rect 11858 8678 11868 8730
rect 11892 8678 11922 8730
rect 11922 8678 11934 8730
rect 11934 8678 11948 8730
rect 11972 8678 11986 8730
rect 11986 8678 11998 8730
rect 11998 8678 12028 8730
rect 12052 8678 12062 8730
rect 12062 8678 12108 8730
rect 11812 8676 11868 8678
rect 11892 8676 11948 8678
rect 11972 8676 12028 8678
rect 12052 8676 12108 8678
rect 17240 8730 17296 8732
rect 17320 8730 17376 8732
rect 17400 8730 17456 8732
rect 17480 8730 17536 8732
rect 17240 8678 17286 8730
rect 17286 8678 17296 8730
rect 17320 8678 17350 8730
rect 17350 8678 17362 8730
rect 17362 8678 17376 8730
rect 17400 8678 17414 8730
rect 17414 8678 17426 8730
rect 17426 8678 17456 8730
rect 17480 8678 17490 8730
rect 17490 8678 17536 8730
rect 17240 8676 17296 8678
rect 17320 8676 17376 8678
rect 17400 8676 17456 8678
rect 17480 8676 17536 8678
rect 3670 8186 3726 8188
rect 3750 8186 3806 8188
rect 3830 8186 3886 8188
rect 3910 8186 3966 8188
rect 3670 8134 3716 8186
rect 3716 8134 3726 8186
rect 3750 8134 3780 8186
rect 3780 8134 3792 8186
rect 3792 8134 3806 8186
rect 3830 8134 3844 8186
rect 3844 8134 3856 8186
rect 3856 8134 3886 8186
rect 3910 8134 3920 8186
rect 3920 8134 3966 8186
rect 3670 8132 3726 8134
rect 3750 8132 3806 8134
rect 3830 8132 3886 8134
rect 3910 8132 3966 8134
rect 9098 8186 9154 8188
rect 9178 8186 9234 8188
rect 9258 8186 9314 8188
rect 9338 8186 9394 8188
rect 9098 8134 9144 8186
rect 9144 8134 9154 8186
rect 9178 8134 9208 8186
rect 9208 8134 9220 8186
rect 9220 8134 9234 8186
rect 9258 8134 9272 8186
rect 9272 8134 9284 8186
rect 9284 8134 9314 8186
rect 9338 8134 9348 8186
rect 9348 8134 9394 8186
rect 9098 8132 9154 8134
rect 9178 8132 9234 8134
rect 9258 8132 9314 8134
rect 9338 8132 9394 8134
rect 14526 8186 14582 8188
rect 14606 8186 14662 8188
rect 14686 8186 14742 8188
rect 14766 8186 14822 8188
rect 14526 8134 14572 8186
rect 14572 8134 14582 8186
rect 14606 8134 14636 8186
rect 14636 8134 14648 8186
rect 14648 8134 14662 8186
rect 14686 8134 14700 8186
rect 14700 8134 14712 8186
rect 14712 8134 14742 8186
rect 14766 8134 14776 8186
rect 14776 8134 14822 8186
rect 14526 8132 14582 8134
rect 14606 8132 14662 8134
rect 14686 8132 14742 8134
rect 14766 8132 14822 8134
rect 19954 21242 20010 21244
rect 20034 21242 20090 21244
rect 20114 21242 20170 21244
rect 20194 21242 20250 21244
rect 19954 21190 20000 21242
rect 20000 21190 20010 21242
rect 20034 21190 20064 21242
rect 20064 21190 20076 21242
rect 20076 21190 20090 21242
rect 20114 21190 20128 21242
rect 20128 21190 20140 21242
rect 20140 21190 20170 21242
rect 20194 21190 20204 21242
rect 20204 21190 20250 21242
rect 19954 21188 20010 21190
rect 20034 21188 20090 21190
rect 20114 21188 20170 21190
rect 20194 21188 20250 21190
rect 19954 20154 20010 20156
rect 20034 20154 20090 20156
rect 20114 20154 20170 20156
rect 20194 20154 20250 20156
rect 19954 20102 20000 20154
rect 20000 20102 20010 20154
rect 20034 20102 20064 20154
rect 20064 20102 20076 20154
rect 20076 20102 20090 20154
rect 20114 20102 20128 20154
rect 20128 20102 20140 20154
rect 20140 20102 20170 20154
rect 20194 20102 20204 20154
rect 20204 20102 20250 20154
rect 19954 20100 20010 20102
rect 20034 20100 20090 20102
rect 20114 20100 20170 20102
rect 20194 20100 20250 20102
rect 19954 19066 20010 19068
rect 20034 19066 20090 19068
rect 20114 19066 20170 19068
rect 20194 19066 20250 19068
rect 19954 19014 20000 19066
rect 20000 19014 20010 19066
rect 20034 19014 20064 19066
rect 20064 19014 20076 19066
rect 20076 19014 20090 19066
rect 20114 19014 20128 19066
rect 20128 19014 20140 19066
rect 20140 19014 20170 19066
rect 20194 19014 20204 19066
rect 20204 19014 20250 19066
rect 19954 19012 20010 19014
rect 20034 19012 20090 19014
rect 20114 19012 20170 19014
rect 20194 19012 20250 19014
rect 19954 17978 20010 17980
rect 20034 17978 20090 17980
rect 20114 17978 20170 17980
rect 20194 17978 20250 17980
rect 19954 17926 20000 17978
rect 20000 17926 20010 17978
rect 20034 17926 20064 17978
rect 20064 17926 20076 17978
rect 20076 17926 20090 17978
rect 20114 17926 20128 17978
rect 20128 17926 20140 17978
rect 20140 17926 20170 17978
rect 20194 17926 20204 17978
rect 20204 17926 20250 17978
rect 19954 17924 20010 17926
rect 20034 17924 20090 17926
rect 20114 17924 20170 17926
rect 20194 17924 20250 17926
rect 19954 16890 20010 16892
rect 20034 16890 20090 16892
rect 20114 16890 20170 16892
rect 20194 16890 20250 16892
rect 19954 16838 20000 16890
rect 20000 16838 20010 16890
rect 20034 16838 20064 16890
rect 20064 16838 20076 16890
rect 20076 16838 20090 16890
rect 20114 16838 20128 16890
rect 20128 16838 20140 16890
rect 20140 16838 20170 16890
rect 20194 16838 20204 16890
rect 20204 16838 20250 16890
rect 19954 16836 20010 16838
rect 20034 16836 20090 16838
rect 20114 16836 20170 16838
rect 20194 16836 20250 16838
rect 19954 15802 20010 15804
rect 20034 15802 20090 15804
rect 20114 15802 20170 15804
rect 20194 15802 20250 15804
rect 19954 15750 20000 15802
rect 20000 15750 20010 15802
rect 20034 15750 20064 15802
rect 20064 15750 20076 15802
rect 20076 15750 20090 15802
rect 20114 15750 20128 15802
rect 20128 15750 20140 15802
rect 20140 15750 20170 15802
rect 20194 15750 20204 15802
rect 20204 15750 20250 15802
rect 19954 15748 20010 15750
rect 20034 15748 20090 15750
rect 20114 15748 20170 15750
rect 20194 15748 20250 15750
rect 19954 14714 20010 14716
rect 20034 14714 20090 14716
rect 20114 14714 20170 14716
rect 20194 14714 20250 14716
rect 19954 14662 20000 14714
rect 20000 14662 20010 14714
rect 20034 14662 20064 14714
rect 20064 14662 20076 14714
rect 20076 14662 20090 14714
rect 20114 14662 20128 14714
rect 20128 14662 20140 14714
rect 20140 14662 20170 14714
rect 20194 14662 20204 14714
rect 20204 14662 20250 14714
rect 19954 14660 20010 14662
rect 20034 14660 20090 14662
rect 20114 14660 20170 14662
rect 20194 14660 20250 14662
rect 19954 13626 20010 13628
rect 20034 13626 20090 13628
rect 20114 13626 20170 13628
rect 20194 13626 20250 13628
rect 19954 13574 20000 13626
rect 20000 13574 20010 13626
rect 20034 13574 20064 13626
rect 20064 13574 20076 13626
rect 20076 13574 20090 13626
rect 20114 13574 20128 13626
rect 20128 13574 20140 13626
rect 20140 13574 20170 13626
rect 20194 13574 20204 13626
rect 20204 13574 20250 13626
rect 19954 13572 20010 13574
rect 20034 13572 20090 13574
rect 20114 13572 20170 13574
rect 20194 13572 20250 13574
rect 22668 20698 22724 20700
rect 22748 20698 22804 20700
rect 22828 20698 22884 20700
rect 22908 20698 22964 20700
rect 22668 20646 22714 20698
rect 22714 20646 22724 20698
rect 22748 20646 22778 20698
rect 22778 20646 22790 20698
rect 22790 20646 22804 20698
rect 22828 20646 22842 20698
rect 22842 20646 22854 20698
rect 22854 20646 22884 20698
rect 22908 20646 22918 20698
rect 22918 20646 22964 20698
rect 22668 20644 22724 20646
rect 22748 20644 22804 20646
rect 22828 20644 22884 20646
rect 22908 20644 22964 20646
rect 22668 19610 22724 19612
rect 22748 19610 22804 19612
rect 22828 19610 22884 19612
rect 22908 19610 22964 19612
rect 22668 19558 22714 19610
rect 22714 19558 22724 19610
rect 22748 19558 22778 19610
rect 22778 19558 22790 19610
rect 22790 19558 22804 19610
rect 22828 19558 22842 19610
rect 22842 19558 22854 19610
rect 22854 19558 22884 19610
rect 22908 19558 22918 19610
rect 22918 19558 22964 19610
rect 22668 19556 22724 19558
rect 22748 19556 22804 19558
rect 22828 19556 22884 19558
rect 22908 19556 22964 19558
rect 22668 18522 22724 18524
rect 22748 18522 22804 18524
rect 22828 18522 22884 18524
rect 22908 18522 22964 18524
rect 22668 18470 22714 18522
rect 22714 18470 22724 18522
rect 22748 18470 22778 18522
rect 22778 18470 22790 18522
rect 22790 18470 22804 18522
rect 22828 18470 22842 18522
rect 22842 18470 22854 18522
rect 22854 18470 22884 18522
rect 22908 18470 22918 18522
rect 22918 18470 22964 18522
rect 22668 18468 22724 18470
rect 22748 18468 22804 18470
rect 22828 18468 22884 18470
rect 22908 18468 22964 18470
rect 22668 17434 22724 17436
rect 22748 17434 22804 17436
rect 22828 17434 22884 17436
rect 22908 17434 22964 17436
rect 22668 17382 22714 17434
rect 22714 17382 22724 17434
rect 22748 17382 22778 17434
rect 22778 17382 22790 17434
rect 22790 17382 22804 17434
rect 22828 17382 22842 17434
rect 22842 17382 22854 17434
rect 22854 17382 22884 17434
rect 22908 17382 22918 17434
rect 22918 17382 22964 17434
rect 22668 17380 22724 17382
rect 22748 17380 22804 17382
rect 22828 17380 22884 17382
rect 22908 17380 22964 17382
rect 22668 16346 22724 16348
rect 22748 16346 22804 16348
rect 22828 16346 22884 16348
rect 22908 16346 22964 16348
rect 22668 16294 22714 16346
rect 22714 16294 22724 16346
rect 22748 16294 22778 16346
rect 22778 16294 22790 16346
rect 22790 16294 22804 16346
rect 22828 16294 22842 16346
rect 22842 16294 22854 16346
rect 22854 16294 22884 16346
rect 22908 16294 22918 16346
rect 22918 16294 22964 16346
rect 22668 16292 22724 16294
rect 22748 16292 22804 16294
rect 22828 16292 22884 16294
rect 22908 16292 22964 16294
rect 22668 15258 22724 15260
rect 22748 15258 22804 15260
rect 22828 15258 22884 15260
rect 22908 15258 22964 15260
rect 22668 15206 22714 15258
rect 22714 15206 22724 15258
rect 22748 15206 22778 15258
rect 22778 15206 22790 15258
rect 22790 15206 22804 15258
rect 22828 15206 22842 15258
rect 22842 15206 22854 15258
rect 22854 15206 22884 15258
rect 22908 15206 22918 15258
rect 22918 15206 22964 15258
rect 22668 15204 22724 15206
rect 22748 15204 22804 15206
rect 22828 15204 22884 15206
rect 22908 15204 22964 15206
rect 22668 14170 22724 14172
rect 22748 14170 22804 14172
rect 22828 14170 22884 14172
rect 22908 14170 22964 14172
rect 22668 14118 22714 14170
rect 22714 14118 22724 14170
rect 22748 14118 22778 14170
rect 22778 14118 22790 14170
rect 22790 14118 22804 14170
rect 22828 14118 22842 14170
rect 22842 14118 22854 14170
rect 22854 14118 22884 14170
rect 22908 14118 22918 14170
rect 22918 14118 22964 14170
rect 22668 14116 22724 14118
rect 22748 14116 22804 14118
rect 22828 14116 22884 14118
rect 22908 14116 22964 14118
rect 22668 13082 22724 13084
rect 22748 13082 22804 13084
rect 22828 13082 22884 13084
rect 22908 13082 22964 13084
rect 22668 13030 22714 13082
rect 22714 13030 22724 13082
rect 22748 13030 22778 13082
rect 22778 13030 22790 13082
rect 22790 13030 22804 13082
rect 22828 13030 22842 13082
rect 22842 13030 22854 13082
rect 22854 13030 22884 13082
rect 22908 13030 22918 13082
rect 22918 13030 22964 13082
rect 22668 13028 22724 13030
rect 22748 13028 22804 13030
rect 22828 13028 22884 13030
rect 22908 13028 22964 13030
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6430 7642
rect 6430 7590 6440 7642
rect 6464 7590 6494 7642
rect 6494 7590 6506 7642
rect 6506 7590 6520 7642
rect 6544 7590 6558 7642
rect 6558 7590 6570 7642
rect 6570 7590 6600 7642
rect 6624 7590 6634 7642
rect 6634 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 11812 7642 11868 7644
rect 11892 7642 11948 7644
rect 11972 7642 12028 7644
rect 12052 7642 12108 7644
rect 11812 7590 11858 7642
rect 11858 7590 11868 7642
rect 11892 7590 11922 7642
rect 11922 7590 11934 7642
rect 11934 7590 11948 7642
rect 11972 7590 11986 7642
rect 11986 7590 11998 7642
rect 11998 7590 12028 7642
rect 12052 7590 12062 7642
rect 12062 7590 12108 7642
rect 11812 7588 11868 7590
rect 11892 7588 11948 7590
rect 11972 7588 12028 7590
rect 12052 7588 12108 7590
rect 17240 7642 17296 7644
rect 17320 7642 17376 7644
rect 17400 7642 17456 7644
rect 17480 7642 17536 7644
rect 17240 7590 17286 7642
rect 17286 7590 17296 7642
rect 17320 7590 17350 7642
rect 17350 7590 17362 7642
rect 17362 7590 17376 7642
rect 17400 7590 17414 7642
rect 17414 7590 17426 7642
rect 17426 7590 17456 7642
rect 17480 7590 17490 7642
rect 17490 7590 17536 7642
rect 17240 7588 17296 7590
rect 17320 7588 17376 7590
rect 17400 7588 17456 7590
rect 17480 7588 17536 7590
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 9098 7098 9154 7100
rect 9178 7098 9234 7100
rect 9258 7098 9314 7100
rect 9338 7098 9394 7100
rect 9098 7046 9144 7098
rect 9144 7046 9154 7098
rect 9178 7046 9208 7098
rect 9208 7046 9220 7098
rect 9220 7046 9234 7098
rect 9258 7046 9272 7098
rect 9272 7046 9284 7098
rect 9284 7046 9314 7098
rect 9338 7046 9348 7098
rect 9348 7046 9394 7098
rect 9098 7044 9154 7046
rect 9178 7044 9234 7046
rect 9258 7044 9314 7046
rect 9338 7044 9394 7046
rect 14526 7098 14582 7100
rect 14606 7098 14662 7100
rect 14686 7098 14742 7100
rect 14766 7098 14822 7100
rect 14526 7046 14572 7098
rect 14572 7046 14582 7098
rect 14606 7046 14636 7098
rect 14636 7046 14648 7098
rect 14648 7046 14662 7098
rect 14686 7046 14700 7098
rect 14700 7046 14712 7098
rect 14712 7046 14742 7098
rect 14766 7046 14776 7098
rect 14776 7046 14822 7098
rect 14526 7044 14582 7046
rect 14606 7044 14662 7046
rect 14686 7044 14742 7046
rect 14766 7044 14822 7046
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6430 6554
rect 6430 6502 6440 6554
rect 6464 6502 6494 6554
rect 6494 6502 6506 6554
rect 6506 6502 6520 6554
rect 6544 6502 6558 6554
rect 6558 6502 6570 6554
rect 6570 6502 6600 6554
rect 6624 6502 6634 6554
rect 6634 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 11812 6554 11868 6556
rect 11892 6554 11948 6556
rect 11972 6554 12028 6556
rect 12052 6554 12108 6556
rect 11812 6502 11858 6554
rect 11858 6502 11868 6554
rect 11892 6502 11922 6554
rect 11922 6502 11934 6554
rect 11934 6502 11948 6554
rect 11972 6502 11986 6554
rect 11986 6502 11998 6554
rect 11998 6502 12028 6554
rect 12052 6502 12062 6554
rect 12062 6502 12108 6554
rect 11812 6500 11868 6502
rect 11892 6500 11948 6502
rect 11972 6500 12028 6502
rect 12052 6500 12108 6502
rect 17240 6554 17296 6556
rect 17320 6554 17376 6556
rect 17400 6554 17456 6556
rect 17480 6554 17536 6556
rect 17240 6502 17286 6554
rect 17286 6502 17296 6554
rect 17320 6502 17350 6554
rect 17350 6502 17362 6554
rect 17362 6502 17376 6554
rect 17400 6502 17414 6554
rect 17414 6502 17426 6554
rect 17426 6502 17456 6554
rect 17480 6502 17490 6554
rect 17490 6502 17536 6554
rect 17240 6500 17296 6502
rect 17320 6500 17376 6502
rect 17400 6500 17456 6502
rect 17480 6500 17536 6502
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 9098 6010 9154 6012
rect 9178 6010 9234 6012
rect 9258 6010 9314 6012
rect 9338 6010 9394 6012
rect 9098 5958 9144 6010
rect 9144 5958 9154 6010
rect 9178 5958 9208 6010
rect 9208 5958 9220 6010
rect 9220 5958 9234 6010
rect 9258 5958 9272 6010
rect 9272 5958 9284 6010
rect 9284 5958 9314 6010
rect 9338 5958 9348 6010
rect 9348 5958 9394 6010
rect 9098 5956 9154 5958
rect 9178 5956 9234 5958
rect 9258 5956 9314 5958
rect 9338 5956 9394 5958
rect 14526 6010 14582 6012
rect 14606 6010 14662 6012
rect 14686 6010 14742 6012
rect 14766 6010 14822 6012
rect 14526 5958 14572 6010
rect 14572 5958 14582 6010
rect 14606 5958 14636 6010
rect 14636 5958 14648 6010
rect 14648 5958 14662 6010
rect 14686 5958 14700 6010
rect 14700 5958 14712 6010
rect 14712 5958 14742 6010
rect 14766 5958 14776 6010
rect 14776 5958 14822 6010
rect 14526 5956 14582 5958
rect 14606 5956 14662 5958
rect 14686 5956 14742 5958
rect 14766 5956 14822 5958
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6430 5466
rect 6430 5414 6440 5466
rect 6464 5414 6494 5466
rect 6494 5414 6506 5466
rect 6506 5414 6520 5466
rect 6544 5414 6558 5466
rect 6558 5414 6570 5466
rect 6570 5414 6600 5466
rect 6624 5414 6634 5466
rect 6634 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 11812 5466 11868 5468
rect 11892 5466 11948 5468
rect 11972 5466 12028 5468
rect 12052 5466 12108 5468
rect 11812 5414 11858 5466
rect 11858 5414 11868 5466
rect 11892 5414 11922 5466
rect 11922 5414 11934 5466
rect 11934 5414 11948 5466
rect 11972 5414 11986 5466
rect 11986 5414 11998 5466
rect 11998 5414 12028 5466
rect 12052 5414 12062 5466
rect 12062 5414 12108 5466
rect 11812 5412 11868 5414
rect 11892 5412 11948 5414
rect 11972 5412 12028 5414
rect 12052 5412 12108 5414
rect 17240 5466 17296 5468
rect 17320 5466 17376 5468
rect 17400 5466 17456 5468
rect 17480 5466 17536 5468
rect 17240 5414 17286 5466
rect 17286 5414 17296 5466
rect 17320 5414 17350 5466
rect 17350 5414 17362 5466
rect 17362 5414 17376 5466
rect 17400 5414 17414 5466
rect 17414 5414 17426 5466
rect 17426 5414 17456 5466
rect 17480 5414 17490 5466
rect 17490 5414 17536 5466
rect 17240 5412 17296 5414
rect 17320 5412 17376 5414
rect 17400 5412 17456 5414
rect 17480 5412 17536 5414
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 9098 4922 9154 4924
rect 9178 4922 9234 4924
rect 9258 4922 9314 4924
rect 9338 4922 9394 4924
rect 9098 4870 9144 4922
rect 9144 4870 9154 4922
rect 9178 4870 9208 4922
rect 9208 4870 9220 4922
rect 9220 4870 9234 4922
rect 9258 4870 9272 4922
rect 9272 4870 9284 4922
rect 9284 4870 9314 4922
rect 9338 4870 9348 4922
rect 9348 4870 9394 4922
rect 9098 4868 9154 4870
rect 9178 4868 9234 4870
rect 9258 4868 9314 4870
rect 9338 4868 9394 4870
rect 14526 4922 14582 4924
rect 14606 4922 14662 4924
rect 14686 4922 14742 4924
rect 14766 4922 14822 4924
rect 14526 4870 14572 4922
rect 14572 4870 14582 4922
rect 14606 4870 14636 4922
rect 14636 4870 14648 4922
rect 14648 4870 14662 4922
rect 14686 4870 14700 4922
rect 14700 4870 14712 4922
rect 14712 4870 14742 4922
rect 14766 4870 14776 4922
rect 14776 4870 14822 4922
rect 14526 4868 14582 4870
rect 14606 4868 14662 4870
rect 14686 4868 14742 4870
rect 14766 4868 14822 4870
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6430 4378
rect 6430 4326 6440 4378
rect 6464 4326 6494 4378
rect 6494 4326 6506 4378
rect 6506 4326 6520 4378
rect 6544 4326 6558 4378
rect 6558 4326 6570 4378
rect 6570 4326 6600 4378
rect 6624 4326 6634 4378
rect 6634 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 11812 4378 11868 4380
rect 11892 4378 11948 4380
rect 11972 4378 12028 4380
rect 12052 4378 12108 4380
rect 11812 4326 11858 4378
rect 11858 4326 11868 4378
rect 11892 4326 11922 4378
rect 11922 4326 11934 4378
rect 11934 4326 11948 4378
rect 11972 4326 11986 4378
rect 11986 4326 11998 4378
rect 11998 4326 12028 4378
rect 12052 4326 12062 4378
rect 12062 4326 12108 4378
rect 11812 4324 11868 4326
rect 11892 4324 11948 4326
rect 11972 4324 12028 4326
rect 12052 4324 12108 4326
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 9098 3834 9154 3836
rect 9178 3834 9234 3836
rect 9258 3834 9314 3836
rect 9338 3834 9394 3836
rect 9098 3782 9144 3834
rect 9144 3782 9154 3834
rect 9178 3782 9208 3834
rect 9208 3782 9220 3834
rect 9220 3782 9234 3834
rect 9258 3782 9272 3834
rect 9272 3782 9284 3834
rect 9284 3782 9314 3834
rect 9338 3782 9348 3834
rect 9348 3782 9394 3834
rect 9098 3780 9154 3782
rect 9178 3780 9234 3782
rect 9258 3780 9314 3782
rect 9338 3780 9394 3782
rect 14526 3834 14582 3836
rect 14606 3834 14662 3836
rect 14686 3834 14742 3836
rect 14766 3834 14822 3836
rect 14526 3782 14572 3834
rect 14572 3782 14582 3834
rect 14606 3782 14636 3834
rect 14636 3782 14648 3834
rect 14648 3782 14662 3834
rect 14686 3782 14700 3834
rect 14700 3782 14712 3834
rect 14712 3782 14742 3834
rect 14766 3782 14776 3834
rect 14776 3782 14822 3834
rect 14526 3780 14582 3782
rect 14606 3780 14662 3782
rect 14686 3780 14742 3782
rect 14766 3780 14822 3782
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6430 3290
rect 6430 3238 6440 3290
rect 6464 3238 6494 3290
rect 6494 3238 6506 3290
rect 6506 3238 6520 3290
rect 6544 3238 6558 3290
rect 6558 3238 6570 3290
rect 6570 3238 6600 3290
rect 6624 3238 6634 3290
rect 6634 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 11812 3290 11868 3292
rect 11892 3290 11948 3292
rect 11972 3290 12028 3292
rect 12052 3290 12108 3292
rect 11812 3238 11858 3290
rect 11858 3238 11868 3290
rect 11892 3238 11922 3290
rect 11922 3238 11934 3290
rect 11934 3238 11948 3290
rect 11972 3238 11986 3290
rect 11986 3238 11998 3290
rect 11998 3238 12028 3290
rect 12052 3238 12062 3290
rect 12062 3238 12108 3290
rect 11812 3236 11868 3238
rect 11892 3236 11948 3238
rect 11972 3236 12028 3238
rect 12052 3236 12108 3238
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 9098 2746 9154 2748
rect 9178 2746 9234 2748
rect 9258 2746 9314 2748
rect 9338 2746 9394 2748
rect 9098 2694 9144 2746
rect 9144 2694 9154 2746
rect 9178 2694 9208 2746
rect 9208 2694 9220 2746
rect 9220 2694 9234 2746
rect 9258 2694 9272 2746
rect 9272 2694 9284 2746
rect 9284 2694 9314 2746
rect 9338 2694 9348 2746
rect 9348 2694 9394 2746
rect 9098 2692 9154 2694
rect 9178 2692 9234 2694
rect 9258 2692 9314 2694
rect 9338 2692 9394 2694
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6430 2202
rect 6430 2150 6440 2202
rect 6464 2150 6494 2202
rect 6494 2150 6506 2202
rect 6506 2150 6520 2202
rect 6544 2150 6558 2202
rect 6558 2150 6570 2202
rect 6570 2150 6600 2202
rect 6624 2150 6634 2202
rect 6634 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 17240 4378 17296 4380
rect 17320 4378 17376 4380
rect 17400 4378 17456 4380
rect 17480 4378 17536 4380
rect 17240 4326 17286 4378
rect 17286 4326 17296 4378
rect 17320 4326 17350 4378
rect 17350 4326 17362 4378
rect 17362 4326 17376 4378
rect 17400 4326 17414 4378
rect 17414 4326 17426 4378
rect 17426 4326 17456 4378
rect 17480 4326 17490 4378
rect 17490 4326 17536 4378
rect 17240 4324 17296 4326
rect 17320 4324 17376 4326
rect 17400 4324 17456 4326
rect 17480 4324 17536 4326
rect 17240 3290 17296 3292
rect 17320 3290 17376 3292
rect 17400 3290 17456 3292
rect 17480 3290 17536 3292
rect 17240 3238 17286 3290
rect 17286 3238 17296 3290
rect 17320 3238 17350 3290
rect 17350 3238 17362 3290
rect 17362 3238 17376 3290
rect 17400 3238 17414 3290
rect 17414 3238 17426 3290
rect 17426 3238 17456 3290
rect 17480 3238 17490 3290
rect 17490 3238 17536 3290
rect 17240 3236 17296 3238
rect 17320 3236 17376 3238
rect 17400 3236 17456 3238
rect 17480 3236 17536 3238
rect 19954 12538 20010 12540
rect 20034 12538 20090 12540
rect 20114 12538 20170 12540
rect 20194 12538 20250 12540
rect 19954 12486 20000 12538
rect 20000 12486 20010 12538
rect 20034 12486 20064 12538
rect 20064 12486 20076 12538
rect 20076 12486 20090 12538
rect 20114 12486 20128 12538
rect 20128 12486 20140 12538
rect 20140 12486 20170 12538
rect 20194 12486 20204 12538
rect 20204 12486 20250 12538
rect 19954 12484 20010 12486
rect 20034 12484 20090 12486
rect 20114 12484 20170 12486
rect 20194 12484 20250 12486
rect 22668 11994 22724 11996
rect 22748 11994 22804 11996
rect 22828 11994 22884 11996
rect 22908 11994 22964 11996
rect 22668 11942 22714 11994
rect 22714 11942 22724 11994
rect 22748 11942 22778 11994
rect 22778 11942 22790 11994
rect 22790 11942 22804 11994
rect 22828 11942 22842 11994
rect 22842 11942 22854 11994
rect 22854 11942 22884 11994
rect 22908 11942 22918 11994
rect 22918 11942 22964 11994
rect 22668 11940 22724 11942
rect 22748 11940 22804 11942
rect 22828 11940 22884 11942
rect 22908 11940 22964 11942
rect 19954 11450 20010 11452
rect 20034 11450 20090 11452
rect 20114 11450 20170 11452
rect 20194 11450 20250 11452
rect 19954 11398 20000 11450
rect 20000 11398 20010 11450
rect 20034 11398 20064 11450
rect 20064 11398 20076 11450
rect 20076 11398 20090 11450
rect 20114 11398 20128 11450
rect 20128 11398 20140 11450
rect 20140 11398 20170 11450
rect 20194 11398 20204 11450
rect 20204 11398 20250 11450
rect 19954 11396 20010 11398
rect 20034 11396 20090 11398
rect 20114 11396 20170 11398
rect 20194 11396 20250 11398
rect 19954 10362 20010 10364
rect 20034 10362 20090 10364
rect 20114 10362 20170 10364
rect 20194 10362 20250 10364
rect 19954 10310 20000 10362
rect 20000 10310 20010 10362
rect 20034 10310 20064 10362
rect 20064 10310 20076 10362
rect 20076 10310 20090 10362
rect 20114 10310 20128 10362
rect 20128 10310 20140 10362
rect 20140 10310 20170 10362
rect 20194 10310 20204 10362
rect 20204 10310 20250 10362
rect 19954 10308 20010 10310
rect 20034 10308 20090 10310
rect 20114 10308 20170 10310
rect 20194 10308 20250 10310
rect 14526 2746 14582 2748
rect 14606 2746 14662 2748
rect 14686 2746 14742 2748
rect 14766 2746 14822 2748
rect 14526 2694 14572 2746
rect 14572 2694 14582 2746
rect 14606 2694 14636 2746
rect 14636 2694 14648 2746
rect 14648 2694 14662 2746
rect 14686 2694 14700 2746
rect 14700 2694 14712 2746
rect 14712 2694 14742 2746
rect 14766 2694 14776 2746
rect 14776 2694 14822 2746
rect 14526 2692 14582 2694
rect 14606 2692 14662 2694
rect 14686 2692 14742 2694
rect 14766 2692 14822 2694
rect 11812 2202 11868 2204
rect 11892 2202 11948 2204
rect 11972 2202 12028 2204
rect 12052 2202 12108 2204
rect 11812 2150 11858 2202
rect 11858 2150 11868 2202
rect 11892 2150 11922 2202
rect 11922 2150 11934 2202
rect 11934 2150 11948 2202
rect 11972 2150 11986 2202
rect 11986 2150 11998 2202
rect 11998 2150 12028 2202
rect 12052 2150 12062 2202
rect 12062 2150 12108 2202
rect 11812 2148 11868 2150
rect 11892 2148 11948 2150
rect 11972 2148 12028 2150
rect 12052 2148 12108 2150
rect 17240 2202 17296 2204
rect 17320 2202 17376 2204
rect 17400 2202 17456 2204
rect 17480 2202 17536 2204
rect 17240 2150 17286 2202
rect 17286 2150 17296 2202
rect 17320 2150 17350 2202
rect 17350 2150 17362 2202
rect 17362 2150 17376 2202
rect 17400 2150 17414 2202
rect 17414 2150 17426 2202
rect 17426 2150 17456 2202
rect 17480 2150 17490 2202
rect 17490 2150 17536 2202
rect 17240 2148 17296 2150
rect 17320 2148 17376 2150
rect 17400 2148 17456 2150
rect 17480 2148 17536 2150
rect 22668 10906 22724 10908
rect 22748 10906 22804 10908
rect 22828 10906 22884 10908
rect 22908 10906 22964 10908
rect 22668 10854 22714 10906
rect 22714 10854 22724 10906
rect 22748 10854 22778 10906
rect 22778 10854 22790 10906
rect 22790 10854 22804 10906
rect 22828 10854 22842 10906
rect 22842 10854 22854 10906
rect 22854 10854 22884 10906
rect 22908 10854 22918 10906
rect 22918 10854 22964 10906
rect 22668 10852 22724 10854
rect 22748 10852 22804 10854
rect 22828 10852 22884 10854
rect 22908 10852 22964 10854
rect 19954 9274 20010 9276
rect 20034 9274 20090 9276
rect 20114 9274 20170 9276
rect 20194 9274 20250 9276
rect 19954 9222 20000 9274
rect 20000 9222 20010 9274
rect 20034 9222 20064 9274
rect 20064 9222 20076 9274
rect 20076 9222 20090 9274
rect 20114 9222 20128 9274
rect 20128 9222 20140 9274
rect 20140 9222 20170 9274
rect 20194 9222 20204 9274
rect 20204 9222 20250 9274
rect 19954 9220 20010 9222
rect 20034 9220 20090 9222
rect 20114 9220 20170 9222
rect 20194 9220 20250 9222
rect 19954 8186 20010 8188
rect 20034 8186 20090 8188
rect 20114 8186 20170 8188
rect 20194 8186 20250 8188
rect 19954 8134 20000 8186
rect 20000 8134 20010 8186
rect 20034 8134 20064 8186
rect 20064 8134 20076 8186
rect 20076 8134 20090 8186
rect 20114 8134 20128 8186
rect 20128 8134 20140 8186
rect 20140 8134 20170 8186
rect 20194 8134 20204 8186
rect 20204 8134 20250 8186
rect 19954 8132 20010 8134
rect 20034 8132 20090 8134
rect 20114 8132 20170 8134
rect 20194 8132 20250 8134
rect 19954 7098 20010 7100
rect 20034 7098 20090 7100
rect 20114 7098 20170 7100
rect 20194 7098 20250 7100
rect 19954 7046 20000 7098
rect 20000 7046 20010 7098
rect 20034 7046 20064 7098
rect 20064 7046 20076 7098
rect 20076 7046 20090 7098
rect 20114 7046 20128 7098
rect 20128 7046 20140 7098
rect 20140 7046 20170 7098
rect 20194 7046 20204 7098
rect 20204 7046 20250 7098
rect 19954 7044 20010 7046
rect 20034 7044 20090 7046
rect 20114 7044 20170 7046
rect 20194 7044 20250 7046
rect 19954 6010 20010 6012
rect 20034 6010 20090 6012
rect 20114 6010 20170 6012
rect 20194 6010 20250 6012
rect 19954 5958 20000 6010
rect 20000 5958 20010 6010
rect 20034 5958 20064 6010
rect 20064 5958 20076 6010
rect 20076 5958 20090 6010
rect 20114 5958 20128 6010
rect 20128 5958 20140 6010
rect 20140 5958 20170 6010
rect 20194 5958 20204 6010
rect 20204 5958 20250 6010
rect 19954 5956 20010 5958
rect 20034 5956 20090 5958
rect 20114 5956 20170 5958
rect 20194 5956 20250 5958
rect 19954 4922 20010 4924
rect 20034 4922 20090 4924
rect 20114 4922 20170 4924
rect 20194 4922 20250 4924
rect 19954 4870 20000 4922
rect 20000 4870 20010 4922
rect 20034 4870 20064 4922
rect 20064 4870 20076 4922
rect 20076 4870 20090 4922
rect 20114 4870 20128 4922
rect 20128 4870 20140 4922
rect 20140 4870 20170 4922
rect 20194 4870 20204 4922
rect 20204 4870 20250 4922
rect 19954 4868 20010 4870
rect 20034 4868 20090 4870
rect 20114 4868 20170 4870
rect 20194 4868 20250 4870
rect 19954 3834 20010 3836
rect 20034 3834 20090 3836
rect 20114 3834 20170 3836
rect 20194 3834 20250 3836
rect 19954 3782 20000 3834
rect 20000 3782 20010 3834
rect 20034 3782 20064 3834
rect 20064 3782 20076 3834
rect 20076 3782 20090 3834
rect 20114 3782 20128 3834
rect 20128 3782 20140 3834
rect 20140 3782 20170 3834
rect 20194 3782 20204 3834
rect 20204 3782 20250 3834
rect 19954 3780 20010 3782
rect 20034 3780 20090 3782
rect 20114 3780 20170 3782
rect 20194 3780 20250 3782
rect 19954 2746 20010 2748
rect 20034 2746 20090 2748
rect 20114 2746 20170 2748
rect 20194 2746 20250 2748
rect 19954 2694 20000 2746
rect 20000 2694 20010 2746
rect 20034 2694 20064 2746
rect 20064 2694 20076 2746
rect 20076 2694 20090 2746
rect 20114 2694 20128 2746
rect 20128 2694 20140 2746
rect 20140 2694 20170 2746
rect 20194 2694 20204 2746
rect 20204 2694 20250 2746
rect 19954 2692 20010 2694
rect 20034 2692 20090 2694
rect 20114 2692 20170 2694
rect 20194 2692 20250 2694
rect 22668 9818 22724 9820
rect 22748 9818 22804 9820
rect 22828 9818 22884 9820
rect 22908 9818 22964 9820
rect 22668 9766 22714 9818
rect 22714 9766 22724 9818
rect 22748 9766 22778 9818
rect 22778 9766 22790 9818
rect 22790 9766 22804 9818
rect 22828 9766 22842 9818
rect 22842 9766 22854 9818
rect 22854 9766 22884 9818
rect 22908 9766 22918 9818
rect 22918 9766 22964 9818
rect 22668 9764 22724 9766
rect 22748 9764 22804 9766
rect 22828 9764 22884 9766
rect 22908 9764 22964 9766
rect 22668 8730 22724 8732
rect 22748 8730 22804 8732
rect 22828 8730 22884 8732
rect 22908 8730 22964 8732
rect 22668 8678 22714 8730
rect 22714 8678 22724 8730
rect 22748 8678 22778 8730
rect 22778 8678 22790 8730
rect 22790 8678 22804 8730
rect 22828 8678 22842 8730
rect 22842 8678 22854 8730
rect 22854 8678 22884 8730
rect 22908 8678 22918 8730
rect 22918 8678 22964 8730
rect 22668 8676 22724 8678
rect 22748 8676 22804 8678
rect 22828 8676 22884 8678
rect 22908 8676 22964 8678
rect 22668 7642 22724 7644
rect 22748 7642 22804 7644
rect 22828 7642 22884 7644
rect 22908 7642 22964 7644
rect 22668 7590 22714 7642
rect 22714 7590 22724 7642
rect 22748 7590 22778 7642
rect 22778 7590 22790 7642
rect 22790 7590 22804 7642
rect 22828 7590 22842 7642
rect 22842 7590 22854 7642
rect 22854 7590 22884 7642
rect 22908 7590 22918 7642
rect 22918 7590 22964 7642
rect 22668 7588 22724 7590
rect 22748 7588 22804 7590
rect 22828 7588 22884 7590
rect 22908 7588 22964 7590
rect 22668 6554 22724 6556
rect 22748 6554 22804 6556
rect 22828 6554 22884 6556
rect 22908 6554 22964 6556
rect 22668 6502 22714 6554
rect 22714 6502 22724 6554
rect 22748 6502 22778 6554
rect 22778 6502 22790 6554
rect 22790 6502 22804 6554
rect 22828 6502 22842 6554
rect 22842 6502 22854 6554
rect 22854 6502 22884 6554
rect 22908 6502 22918 6554
rect 22918 6502 22964 6554
rect 22668 6500 22724 6502
rect 22748 6500 22804 6502
rect 22828 6500 22884 6502
rect 22908 6500 22964 6502
rect 22668 5466 22724 5468
rect 22748 5466 22804 5468
rect 22828 5466 22884 5468
rect 22908 5466 22964 5468
rect 22668 5414 22714 5466
rect 22714 5414 22724 5466
rect 22748 5414 22778 5466
rect 22778 5414 22790 5466
rect 22790 5414 22804 5466
rect 22828 5414 22842 5466
rect 22842 5414 22854 5466
rect 22854 5414 22884 5466
rect 22908 5414 22918 5466
rect 22918 5414 22964 5466
rect 22668 5412 22724 5414
rect 22748 5412 22804 5414
rect 22828 5412 22884 5414
rect 22908 5412 22964 5414
rect 22668 4378 22724 4380
rect 22748 4378 22804 4380
rect 22828 4378 22884 4380
rect 22908 4378 22964 4380
rect 22668 4326 22714 4378
rect 22714 4326 22724 4378
rect 22748 4326 22778 4378
rect 22778 4326 22790 4378
rect 22790 4326 22804 4378
rect 22828 4326 22842 4378
rect 22842 4326 22854 4378
rect 22854 4326 22884 4378
rect 22908 4326 22918 4378
rect 22918 4326 22964 4378
rect 22668 4324 22724 4326
rect 22748 4324 22804 4326
rect 22828 4324 22884 4326
rect 22908 4324 22964 4326
rect 22668 3290 22724 3292
rect 22748 3290 22804 3292
rect 22828 3290 22884 3292
rect 22908 3290 22964 3292
rect 22668 3238 22714 3290
rect 22714 3238 22724 3290
rect 22748 3238 22778 3290
rect 22778 3238 22790 3290
rect 22790 3238 22804 3290
rect 22828 3238 22842 3290
rect 22842 3238 22854 3290
rect 22854 3238 22884 3290
rect 22908 3238 22918 3290
rect 22918 3238 22964 3290
rect 22668 3236 22724 3238
rect 22748 3236 22804 3238
rect 22828 3236 22884 3238
rect 22908 3236 22964 3238
rect 22668 2202 22724 2204
rect 22748 2202 22804 2204
rect 22828 2202 22884 2204
rect 22908 2202 22964 2204
rect 22668 2150 22714 2202
rect 22714 2150 22724 2202
rect 22748 2150 22778 2202
rect 22778 2150 22790 2202
rect 22790 2150 22804 2202
rect 22828 2150 22842 2202
rect 22842 2150 22854 2202
rect 22854 2150 22884 2202
rect 22908 2150 22918 2202
rect 22918 2150 22964 2202
rect 22668 2148 22724 2150
rect 22748 2148 22804 2150
rect 22828 2148 22884 2150
rect 22908 2148 22964 2150
<< metal3 >>
rect 6374 21792 6690 21793
rect 6374 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6690 21792
rect 6374 21727 6690 21728
rect 11802 21792 12118 21793
rect 11802 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12118 21792
rect 11802 21727 12118 21728
rect 17230 21792 17546 21793
rect 17230 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17546 21792
rect 17230 21727 17546 21728
rect 22658 21792 22974 21793
rect 22658 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22974 21792
rect 22658 21727 22974 21728
rect 3660 21248 3976 21249
rect 3660 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3976 21248
rect 3660 21183 3976 21184
rect 9088 21248 9404 21249
rect 9088 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9404 21248
rect 9088 21183 9404 21184
rect 14516 21248 14832 21249
rect 14516 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14832 21248
rect 14516 21183 14832 21184
rect 19944 21248 20260 21249
rect 19944 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20260 21248
rect 19944 21183 20260 21184
rect 6374 20704 6690 20705
rect 6374 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6690 20704
rect 6374 20639 6690 20640
rect 11802 20704 12118 20705
rect 11802 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12118 20704
rect 11802 20639 12118 20640
rect 17230 20704 17546 20705
rect 17230 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17546 20704
rect 17230 20639 17546 20640
rect 22658 20704 22974 20705
rect 22658 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22974 20704
rect 22658 20639 22974 20640
rect 3660 20160 3976 20161
rect 3660 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3976 20160
rect 3660 20095 3976 20096
rect 9088 20160 9404 20161
rect 9088 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9404 20160
rect 9088 20095 9404 20096
rect 14516 20160 14832 20161
rect 14516 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14832 20160
rect 14516 20095 14832 20096
rect 19944 20160 20260 20161
rect 19944 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20260 20160
rect 19944 20095 20260 20096
rect 6374 19616 6690 19617
rect 6374 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6690 19616
rect 6374 19551 6690 19552
rect 11802 19616 12118 19617
rect 11802 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12118 19616
rect 11802 19551 12118 19552
rect 17230 19616 17546 19617
rect 17230 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17546 19616
rect 17230 19551 17546 19552
rect 22658 19616 22974 19617
rect 22658 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22974 19616
rect 22658 19551 22974 19552
rect 3660 19072 3976 19073
rect 3660 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3976 19072
rect 3660 19007 3976 19008
rect 9088 19072 9404 19073
rect 9088 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9404 19072
rect 9088 19007 9404 19008
rect 14516 19072 14832 19073
rect 14516 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14832 19072
rect 14516 19007 14832 19008
rect 19944 19072 20260 19073
rect 19944 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20260 19072
rect 19944 19007 20260 19008
rect 6374 18528 6690 18529
rect 6374 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6690 18528
rect 6374 18463 6690 18464
rect 11802 18528 12118 18529
rect 11802 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12118 18528
rect 11802 18463 12118 18464
rect 17230 18528 17546 18529
rect 17230 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17546 18528
rect 17230 18463 17546 18464
rect 22658 18528 22974 18529
rect 22658 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22974 18528
rect 22658 18463 22974 18464
rect 3660 17984 3976 17985
rect 3660 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3976 17984
rect 3660 17919 3976 17920
rect 9088 17984 9404 17985
rect 9088 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9404 17984
rect 9088 17919 9404 17920
rect 14516 17984 14832 17985
rect 14516 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14832 17984
rect 14516 17919 14832 17920
rect 19944 17984 20260 17985
rect 19944 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20260 17984
rect 19944 17919 20260 17920
rect 6374 17440 6690 17441
rect 6374 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6690 17440
rect 6374 17375 6690 17376
rect 11802 17440 12118 17441
rect 11802 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12118 17440
rect 11802 17375 12118 17376
rect 17230 17440 17546 17441
rect 17230 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17546 17440
rect 17230 17375 17546 17376
rect 22658 17440 22974 17441
rect 22658 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22974 17440
rect 22658 17375 22974 17376
rect 3660 16896 3976 16897
rect 3660 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3976 16896
rect 3660 16831 3976 16832
rect 9088 16896 9404 16897
rect 9088 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9404 16896
rect 9088 16831 9404 16832
rect 14516 16896 14832 16897
rect 14516 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14832 16896
rect 14516 16831 14832 16832
rect 19944 16896 20260 16897
rect 19944 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20260 16896
rect 19944 16831 20260 16832
rect 6374 16352 6690 16353
rect 6374 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6690 16352
rect 6374 16287 6690 16288
rect 11802 16352 12118 16353
rect 11802 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12118 16352
rect 11802 16287 12118 16288
rect 17230 16352 17546 16353
rect 17230 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17546 16352
rect 17230 16287 17546 16288
rect 22658 16352 22974 16353
rect 22658 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22974 16352
rect 22658 16287 22974 16288
rect 3660 15808 3976 15809
rect 3660 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3976 15808
rect 3660 15743 3976 15744
rect 9088 15808 9404 15809
rect 9088 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9404 15808
rect 9088 15743 9404 15744
rect 14516 15808 14832 15809
rect 14516 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14832 15808
rect 14516 15743 14832 15744
rect 19944 15808 20260 15809
rect 19944 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20260 15808
rect 19944 15743 20260 15744
rect 6374 15264 6690 15265
rect 6374 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6690 15264
rect 6374 15199 6690 15200
rect 11802 15264 12118 15265
rect 11802 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12118 15264
rect 11802 15199 12118 15200
rect 17230 15264 17546 15265
rect 17230 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17546 15264
rect 17230 15199 17546 15200
rect 22658 15264 22974 15265
rect 22658 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22974 15264
rect 22658 15199 22974 15200
rect 3660 14720 3976 14721
rect 3660 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3976 14720
rect 3660 14655 3976 14656
rect 9088 14720 9404 14721
rect 9088 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9404 14720
rect 9088 14655 9404 14656
rect 14516 14720 14832 14721
rect 14516 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14832 14720
rect 14516 14655 14832 14656
rect 19944 14720 20260 14721
rect 19944 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20260 14720
rect 19944 14655 20260 14656
rect 6374 14176 6690 14177
rect 6374 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6690 14176
rect 6374 14111 6690 14112
rect 11802 14176 12118 14177
rect 11802 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12118 14176
rect 11802 14111 12118 14112
rect 17230 14176 17546 14177
rect 17230 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17546 14176
rect 17230 14111 17546 14112
rect 22658 14176 22974 14177
rect 22658 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22974 14176
rect 22658 14111 22974 14112
rect 3660 13632 3976 13633
rect 3660 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3976 13632
rect 3660 13567 3976 13568
rect 9088 13632 9404 13633
rect 9088 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9404 13632
rect 9088 13567 9404 13568
rect 14516 13632 14832 13633
rect 14516 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14832 13632
rect 14516 13567 14832 13568
rect 19944 13632 20260 13633
rect 19944 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20260 13632
rect 19944 13567 20260 13568
rect 6374 13088 6690 13089
rect 6374 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6690 13088
rect 6374 13023 6690 13024
rect 11802 13088 12118 13089
rect 11802 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12118 13088
rect 11802 13023 12118 13024
rect 17230 13088 17546 13089
rect 17230 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17546 13088
rect 17230 13023 17546 13024
rect 22658 13088 22974 13089
rect 22658 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22974 13088
rect 22658 13023 22974 13024
rect 3660 12544 3976 12545
rect 3660 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3976 12544
rect 3660 12479 3976 12480
rect 9088 12544 9404 12545
rect 9088 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9404 12544
rect 9088 12479 9404 12480
rect 14516 12544 14832 12545
rect 14516 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14832 12544
rect 14516 12479 14832 12480
rect 19944 12544 20260 12545
rect 19944 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20260 12544
rect 19944 12479 20260 12480
rect 6374 12000 6690 12001
rect 6374 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6690 12000
rect 6374 11935 6690 11936
rect 11802 12000 12118 12001
rect 11802 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12118 12000
rect 11802 11935 12118 11936
rect 17230 12000 17546 12001
rect 17230 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17546 12000
rect 17230 11935 17546 11936
rect 22658 12000 22974 12001
rect 22658 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22974 12000
rect 22658 11935 22974 11936
rect 3660 11456 3976 11457
rect 3660 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3976 11456
rect 3660 11391 3976 11392
rect 9088 11456 9404 11457
rect 9088 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9404 11456
rect 9088 11391 9404 11392
rect 14516 11456 14832 11457
rect 14516 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14832 11456
rect 14516 11391 14832 11392
rect 19944 11456 20260 11457
rect 19944 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20260 11456
rect 19944 11391 20260 11392
rect 6374 10912 6690 10913
rect 6374 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6690 10912
rect 6374 10847 6690 10848
rect 11802 10912 12118 10913
rect 11802 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12118 10912
rect 11802 10847 12118 10848
rect 17230 10912 17546 10913
rect 17230 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17546 10912
rect 17230 10847 17546 10848
rect 22658 10912 22974 10913
rect 22658 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22974 10912
rect 22658 10847 22974 10848
rect 3660 10368 3976 10369
rect 3660 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3976 10368
rect 3660 10303 3976 10304
rect 9088 10368 9404 10369
rect 9088 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9404 10368
rect 9088 10303 9404 10304
rect 14516 10368 14832 10369
rect 14516 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14832 10368
rect 14516 10303 14832 10304
rect 19944 10368 20260 10369
rect 19944 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20260 10368
rect 19944 10303 20260 10304
rect 6374 9824 6690 9825
rect 6374 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6690 9824
rect 6374 9759 6690 9760
rect 11802 9824 12118 9825
rect 11802 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12118 9824
rect 11802 9759 12118 9760
rect 17230 9824 17546 9825
rect 17230 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17546 9824
rect 17230 9759 17546 9760
rect 22658 9824 22974 9825
rect 22658 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22974 9824
rect 22658 9759 22974 9760
rect 3660 9280 3976 9281
rect 3660 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3976 9280
rect 3660 9215 3976 9216
rect 9088 9280 9404 9281
rect 9088 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9404 9280
rect 9088 9215 9404 9216
rect 14516 9280 14832 9281
rect 14516 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14832 9280
rect 14516 9215 14832 9216
rect 19944 9280 20260 9281
rect 19944 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20260 9280
rect 19944 9215 20260 9216
rect 6374 8736 6690 8737
rect 6374 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6690 8736
rect 6374 8671 6690 8672
rect 11802 8736 12118 8737
rect 11802 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12118 8736
rect 11802 8671 12118 8672
rect 17230 8736 17546 8737
rect 17230 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17546 8736
rect 17230 8671 17546 8672
rect 22658 8736 22974 8737
rect 22658 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22974 8736
rect 22658 8671 22974 8672
rect 3660 8192 3976 8193
rect 3660 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3976 8192
rect 3660 8127 3976 8128
rect 9088 8192 9404 8193
rect 9088 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9404 8192
rect 9088 8127 9404 8128
rect 14516 8192 14832 8193
rect 14516 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14832 8192
rect 14516 8127 14832 8128
rect 19944 8192 20260 8193
rect 19944 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20260 8192
rect 19944 8127 20260 8128
rect 6374 7648 6690 7649
rect 6374 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6690 7648
rect 6374 7583 6690 7584
rect 11802 7648 12118 7649
rect 11802 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12118 7648
rect 11802 7583 12118 7584
rect 17230 7648 17546 7649
rect 17230 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17546 7648
rect 17230 7583 17546 7584
rect 22658 7648 22974 7649
rect 22658 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22974 7648
rect 22658 7583 22974 7584
rect 3660 7104 3976 7105
rect 3660 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3976 7104
rect 3660 7039 3976 7040
rect 9088 7104 9404 7105
rect 9088 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9404 7104
rect 9088 7039 9404 7040
rect 14516 7104 14832 7105
rect 14516 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14832 7104
rect 14516 7039 14832 7040
rect 19944 7104 20260 7105
rect 19944 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20260 7104
rect 19944 7039 20260 7040
rect 6374 6560 6690 6561
rect 6374 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6690 6560
rect 6374 6495 6690 6496
rect 11802 6560 12118 6561
rect 11802 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12118 6560
rect 11802 6495 12118 6496
rect 17230 6560 17546 6561
rect 17230 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17546 6560
rect 17230 6495 17546 6496
rect 22658 6560 22974 6561
rect 22658 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22974 6560
rect 22658 6495 22974 6496
rect 3660 6016 3976 6017
rect 3660 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3976 6016
rect 3660 5951 3976 5952
rect 9088 6016 9404 6017
rect 9088 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9404 6016
rect 9088 5951 9404 5952
rect 14516 6016 14832 6017
rect 14516 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14832 6016
rect 14516 5951 14832 5952
rect 19944 6016 20260 6017
rect 19944 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20260 6016
rect 19944 5951 20260 5952
rect 6374 5472 6690 5473
rect 6374 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6690 5472
rect 6374 5407 6690 5408
rect 11802 5472 12118 5473
rect 11802 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12118 5472
rect 11802 5407 12118 5408
rect 17230 5472 17546 5473
rect 17230 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17546 5472
rect 17230 5407 17546 5408
rect 22658 5472 22974 5473
rect 22658 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22974 5472
rect 22658 5407 22974 5408
rect 3660 4928 3976 4929
rect 3660 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3976 4928
rect 3660 4863 3976 4864
rect 9088 4928 9404 4929
rect 9088 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9404 4928
rect 9088 4863 9404 4864
rect 14516 4928 14832 4929
rect 14516 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14832 4928
rect 14516 4863 14832 4864
rect 19944 4928 20260 4929
rect 19944 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20260 4928
rect 19944 4863 20260 4864
rect 6374 4384 6690 4385
rect 6374 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6690 4384
rect 6374 4319 6690 4320
rect 11802 4384 12118 4385
rect 11802 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12118 4384
rect 11802 4319 12118 4320
rect 17230 4384 17546 4385
rect 17230 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17546 4384
rect 17230 4319 17546 4320
rect 22658 4384 22974 4385
rect 22658 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22974 4384
rect 22658 4319 22974 4320
rect 3660 3840 3976 3841
rect 3660 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3976 3840
rect 3660 3775 3976 3776
rect 9088 3840 9404 3841
rect 9088 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9404 3840
rect 9088 3775 9404 3776
rect 14516 3840 14832 3841
rect 14516 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14832 3840
rect 14516 3775 14832 3776
rect 19944 3840 20260 3841
rect 19944 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20260 3840
rect 19944 3775 20260 3776
rect 6374 3296 6690 3297
rect 6374 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6690 3296
rect 6374 3231 6690 3232
rect 11802 3296 12118 3297
rect 11802 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12118 3296
rect 11802 3231 12118 3232
rect 17230 3296 17546 3297
rect 17230 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17546 3296
rect 17230 3231 17546 3232
rect 22658 3296 22974 3297
rect 22658 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22974 3296
rect 22658 3231 22974 3232
rect 3660 2752 3976 2753
rect 3660 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3976 2752
rect 3660 2687 3976 2688
rect 9088 2752 9404 2753
rect 9088 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9404 2752
rect 9088 2687 9404 2688
rect 14516 2752 14832 2753
rect 14516 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14832 2752
rect 14516 2687 14832 2688
rect 19944 2752 20260 2753
rect 19944 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20260 2752
rect 19944 2687 20260 2688
rect 6374 2208 6690 2209
rect 6374 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6690 2208
rect 6374 2143 6690 2144
rect 11802 2208 12118 2209
rect 11802 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12118 2208
rect 11802 2143 12118 2144
rect 17230 2208 17546 2209
rect 17230 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17546 2208
rect 17230 2143 17546 2144
rect 22658 2208 22974 2209
rect 22658 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22974 2208
rect 22658 2143 22974 2144
<< via3 >>
rect 6380 21788 6444 21792
rect 6380 21732 6384 21788
rect 6384 21732 6440 21788
rect 6440 21732 6444 21788
rect 6380 21728 6444 21732
rect 6460 21788 6524 21792
rect 6460 21732 6464 21788
rect 6464 21732 6520 21788
rect 6520 21732 6524 21788
rect 6460 21728 6524 21732
rect 6540 21788 6604 21792
rect 6540 21732 6544 21788
rect 6544 21732 6600 21788
rect 6600 21732 6604 21788
rect 6540 21728 6604 21732
rect 6620 21788 6684 21792
rect 6620 21732 6624 21788
rect 6624 21732 6680 21788
rect 6680 21732 6684 21788
rect 6620 21728 6684 21732
rect 11808 21788 11872 21792
rect 11808 21732 11812 21788
rect 11812 21732 11868 21788
rect 11868 21732 11872 21788
rect 11808 21728 11872 21732
rect 11888 21788 11952 21792
rect 11888 21732 11892 21788
rect 11892 21732 11948 21788
rect 11948 21732 11952 21788
rect 11888 21728 11952 21732
rect 11968 21788 12032 21792
rect 11968 21732 11972 21788
rect 11972 21732 12028 21788
rect 12028 21732 12032 21788
rect 11968 21728 12032 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 17316 21788 17380 21792
rect 17316 21732 17320 21788
rect 17320 21732 17376 21788
rect 17376 21732 17380 21788
rect 17316 21728 17380 21732
rect 17396 21788 17460 21792
rect 17396 21732 17400 21788
rect 17400 21732 17456 21788
rect 17456 21732 17460 21788
rect 17396 21728 17460 21732
rect 17476 21788 17540 21792
rect 17476 21732 17480 21788
rect 17480 21732 17536 21788
rect 17536 21732 17540 21788
rect 17476 21728 17540 21732
rect 22664 21788 22728 21792
rect 22664 21732 22668 21788
rect 22668 21732 22724 21788
rect 22724 21732 22728 21788
rect 22664 21728 22728 21732
rect 22744 21788 22808 21792
rect 22744 21732 22748 21788
rect 22748 21732 22804 21788
rect 22804 21732 22808 21788
rect 22744 21728 22808 21732
rect 22824 21788 22888 21792
rect 22824 21732 22828 21788
rect 22828 21732 22884 21788
rect 22884 21732 22888 21788
rect 22824 21728 22888 21732
rect 22904 21788 22968 21792
rect 22904 21732 22908 21788
rect 22908 21732 22964 21788
rect 22964 21732 22968 21788
rect 22904 21728 22968 21732
rect 3666 21244 3730 21248
rect 3666 21188 3670 21244
rect 3670 21188 3726 21244
rect 3726 21188 3730 21244
rect 3666 21184 3730 21188
rect 3746 21244 3810 21248
rect 3746 21188 3750 21244
rect 3750 21188 3806 21244
rect 3806 21188 3810 21244
rect 3746 21184 3810 21188
rect 3826 21244 3890 21248
rect 3826 21188 3830 21244
rect 3830 21188 3886 21244
rect 3886 21188 3890 21244
rect 3826 21184 3890 21188
rect 3906 21244 3970 21248
rect 3906 21188 3910 21244
rect 3910 21188 3966 21244
rect 3966 21188 3970 21244
rect 3906 21184 3970 21188
rect 9094 21244 9158 21248
rect 9094 21188 9098 21244
rect 9098 21188 9154 21244
rect 9154 21188 9158 21244
rect 9094 21184 9158 21188
rect 9174 21244 9238 21248
rect 9174 21188 9178 21244
rect 9178 21188 9234 21244
rect 9234 21188 9238 21244
rect 9174 21184 9238 21188
rect 9254 21244 9318 21248
rect 9254 21188 9258 21244
rect 9258 21188 9314 21244
rect 9314 21188 9318 21244
rect 9254 21184 9318 21188
rect 9334 21244 9398 21248
rect 9334 21188 9338 21244
rect 9338 21188 9394 21244
rect 9394 21188 9398 21244
rect 9334 21184 9398 21188
rect 14522 21244 14586 21248
rect 14522 21188 14526 21244
rect 14526 21188 14582 21244
rect 14582 21188 14586 21244
rect 14522 21184 14586 21188
rect 14602 21244 14666 21248
rect 14602 21188 14606 21244
rect 14606 21188 14662 21244
rect 14662 21188 14666 21244
rect 14602 21184 14666 21188
rect 14682 21244 14746 21248
rect 14682 21188 14686 21244
rect 14686 21188 14742 21244
rect 14742 21188 14746 21244
rect 14682 21184 14746 21188
rect 14762 21244 14826 21248
rect 14762 21188 14766 21244
rect 14766 21188 14822 21244
rect 14822 21188 14826 21244
rect 14762 21184 14826 21188
rect 19950 21244 20014 21248
rect 19950 21188 19954 21244
rect 19954 21188 20010 21244
rect 20010 21188 20014 21244
rect 19950 21184 20014 21188
rect 20030 21244 20094 21248
rect 20030 21188 20034 21244
rect 20034 21188 20090 21244
rect 20090 21188 20094 21244
rect 20030 21184 20094 21188
rect 20110 21244 20174 21248
rect 20110 21188 20114 21244
rect 20114 21188 20170 21244
rect 20170 21188 20174 21244
rect 20110 21184 20174 21188
rect 20190 21244 20254 21248
rect 20190 21188 20194 21244
rect 20194 21188 20250 21244
rect 20250 21188 20254 21244
rect 20190 21184 20254 21188
rect 6380 20700 6444 20704
rect 6380 20644 6384 20700
rect 6384 20644 6440 20700
rect 6440 20644 6444 20700
rect 6380 20640 6444 20644
rect 6460 20700 6524 20704
rect 6460 20644 6464 20700
rect 6464 20644 6520 20700
rect 6520 20644 6524 20700
rect 6460 20640 6524 20644
rect 6540 20700 6604 20704
rect 6540 20644 6544 20700
rect 6544 20644 6600 20700
rect 6600 20644 6604 20700
rect 6540 20640 6604 20644
rect 6620 20700 6684 20704
rect 6620 20644 6624 20700
rect 6624 20644 6680 20700
rect 6680 20644 6684 20700
rect 6620 20640 6684 20644
rect 11808 20700 11872 20704
rect 11808 20644 11812 20700
rect 11812 20644 11868 20700
rect 11868 20644 11872 20700
rect 11808 20640 11872 20644
rect 11888 20700 11952 20704
rect 11888 20644 11892 20700
rect 11892 20644 11948 20700
rect 11948 20644 11952 20700
rect 11888 20640 11952 20644
rect 11968 20700 12032 20704
rect 11968 20644 11972 20700
rect 11972 20644 12028 20700
rect 12028 20644 12032 20700
rect 11968 20640 12032 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 17316 20700 17380 20704
rect 17316 20644 17320 20700
rect 17320 20644 17376 20700
rect 17376 20644 17380 20700
rect 17316 20640 17380 20644
rect 17396 20700 17460 20704
rect 17396 20644 17400 20700
rect 17400 20644 17456 20700
rect 17456 20644 17460 20700
rect 17396 20640 17460 20644
rect 17476 20700 17540 20704
rect 17476 20644 17480 20700
rect 17480 20644 17536 20700
rect 17536 20644 17540 20700
rect 17476 20640 17540 20644
rect 22664 20700 22728 20704
rect 22664 20644 22668 20700
rect 22668 20644 22724 20700
rect 22724 20644 22728 20700
rect 22664 20640 22728 20644
rect 22744 20700 22808 20704
rect 22744 20644 22748 20700
rect 22748 20644 22804 20700
rect 22804 20644 22808 20700
rect 22744 20640 22808 20644
rect 22824 20700 22888 20704
rect 22824 20644 22828 20700
rect 22828 20644 22884 20700
rect 22884 20644 22888 20700
rect 22824 20640 22888 20644
rect 22904 20700 22968 20704
rect 22904 20644 22908 20700
rect 22908 20644 22964 20700
rect 22964 20644 22968 20700
rect 22904 20640 22968 20644
rect 3666 20156 3730 20160
rect 3666 20100 3670 20156
rect 3670 20100 3726 20156
rect 3726 20100 3730 20156
rect 3666 20096 3730 20100
rect 3746 20156 3810 20160
rect 3746 20100 3750 20156
rect 3750 20100 3806 20156
rect 3806 20100 3810 20156
rect 3746 20096 3810 20100
rect 3826 20156 3890 20160
rect 3826 20100 3830 20156
rect 3830 20100 3886 20156
rect 3886 20100 3890 20156
rect 3826 20096 3890 20100
rect 3906 20156 3970 20160
rect 3906 20100 3910 20156
rect 3910 20100 3966 20156
rect 3966 20100 3970 20156
rect 3906 20096 3970 20100
rect 9094 20156 9158 20160
rect 9094 20100 9098 20156
rect 9098 20100 9154 20156
rect 9154 20100 9158 20156
rect 9094 20096 9158 20100
rect 9174 20156 9238 20160
rect 9174 20100 9178 20156
rect 9178 20100 9234 20156
rect 9234 20100 9238 20156
rect 9174 20096 9238 20100
rect 9254 20156 9318 20160
rect 9254 20100 9258 20156
rect 9258 20100 9314 20156
rect 9314 20100 9318 20156
rect 9254 20096 9318 20100
rect 9334 20156 9398 20160
rect 9334 20100 9338 20156
rect 9338 20100 9394 20156
rect 9394 20100 9398 20156
rect 9334 20096 9398 20100
rect 14522 20156 14586 20160
rect 14522 20100 14526 20156
rect 14526 20100 14582 20156
rect 14582 20100 14586 20156
rect 14522 20096 14586 20100
rect 14602 20156 14666 20160
rect 14602 20100 14606 20156
rect 14606 20100 14662 20156
rect 14662 20100 14666 20156
rect 14602 20096 14666 20100
rect 14682 20156 14746 20160
rect 14682 20100 14686 20156
rect 14686 20100 14742 20156
rect 14742 20100 14746 20156
rect 14682 20096 14746 20100
rect 14762 20156 14826 20160
rect 14762 20100 14766 20156
rect 14766 20100 14822 20156
rect 14822 20100 14826 20156
rect 14762 20096 14826 20100
rect 19950 20156 20014 20160
rect 19950 20100 19954 20156
rect 19954 20100 20010 20156
rect 20010 20100 20014 20156
rect 19950 20096 20014 20100
rect 20030 20156 20094 20160
rect 20030 20100 20034 20156
rect 20034 20100 20090 20156
rect 20090 20100 20094 20156
rect 20030 20096 20094 20100
rect 20110 20156 20174 20160
rect 20110 20100 20114 20156
rect 20114 20100 20170 20156
rect 20170 20100 20174 20156
rect 20110 20096 20174 20100
rect 20190 20156 20254 20160
rect 20190 20100 20194 20156
rect 20194 20100 20250 20156
rect 20250 20100 20254 20156
rect 20190 20096 20254 20100
rect 6380 19612 6444 19616
rect 6380 19556 6384 19612
rect 6384 19556 6440 19612
rect 6440 19556 6444 19612
rect 6380 19552 6444 19556
rect 6460 19612 6524 19616
rect 6460 19556 6464 19612
rect 6464 19556 6520 19612
rect 6520 19556 6524 19612
rect 6460 19552 6524 19556
rect 6540 19612 6604 19616
rect 6540 19556 6544 19612
rect 6544 19556 6600 19612
rect 6600 19556 6604 19612
rect 6540 19552 6604 19556
rect 6620 19612 6684 19616
rect 6620 19556 6624 19612
rect 6624 19556 6680 19612
rect 6680 19556 6684 19612
rect 6620 19552 6684 19556
rect 11808 19612 11872 19616
rect 11808 19556 11812 19612
rect 11812 19556 11868 19612
rect 11868 19556 11872 19612
rect 11808 19552 11872 19556
rect 11888 19612 11952 19616
rect 11888 19556 11892 19612
rect 11892 19556 11948 19612
rect 11948 19556 11952 19612
rect 11888 19552 11952 19556
rect 11968 19612 12032 19616
rect 11968 19556 11972 19612
rect 11972 19556 12028 19612
rect 12028 19556 12032 19612
rect 11968 19552 12032 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 17316 19612 17380 19616
rect 17316 19556 17320 19612
rect 17320 19556 17376 19612
rect 17376 19556 17380 19612
rect 17316 19552 17380 19556
rect 17396 19612 17460 19616
rect 17396 19556 17400 19612
rect 17400 19556 17456 19612
rect 17456 19556 17460 19612
rect 17396 19552 17460 19556
rect 17476 19612 17540 19616
rect 17476 19556 17480 19612
rect 17480 19556 17536 19612
rect 17536 19556 17540 19612
rect 17476 19552 17540 19556
rect 22664 19612 22728 19616
rect 22664 19556 22668 19612
rect 22668 19556 22724 19612
rect 22724 19556 22728 19612
rect 22664 19552 22728 19556
rect 22744 19612 22808 19616
rect 22744 19556 22748 19612
rect 22748 19556 22804 19612
rect 22804 19556 22808 19612
rect 22744 19552 22808 19556
rect 22824 19612 22888 19616
rect 22824 19556 22828 19612
rect 22828 19556 22884 19612
rect 22884 19556 22888 19612
rect 22824 19552 22888 19556
rect 22904 19612 22968 19616
rect 22904 19556 22908 19612
rect 22908 19556 22964 19612
rect 22964 19556 22968 19612
rect 22904 19552 22968 19556
rect 3666 19068 3730 19072
rect 3666 19012 3670 19068
rect 3670 19012 3726 19068
rect 3726 19012 3730 19068
rect 3666 19008 3730 19012
rect 3746 19068 3810 19072
rect 3746 19012 3750 19068
rect 3750 19012 3806 19068
rect 3806 19012 3810 19068
rect 3746 19008 3810 19012
rect 3826 19068 3890 19072
rect 3826 19012 3830 19068
rect 3830 19012 3886 19068
rect 3886 19012 3890 19068
rect 3826 19008 3890 19012
rect 3906 19068 3970 19072
rect 3906 19012 3910 19068
rect 3910 19012 3966 19068
rect 3966 19012 3970 19068
rect 3906 19008 3970 19012
rect 9094 19068 9158 19072
rect 9094 19012 9098 19068
rect 9098 19012 9154 19068
rect 9154 19012 9158 19068
rect 9094 19008 9158 19012
rect 9174 19068 9238 19072
rect 9174 19012 9178 19068
rect 9178 19012 9234 19068
rect 9234 19012 9238 19068
rect 9174 19008 9238 19012
rect 9254 19068 9318 19072
rect 9254 19012 9258 19068
rect 9258 19012 9314 19068
rect 9314 19012 9318 19068
rect 9254 19008 9318 19012
rect 9334 19068 9398 19072
rect 9334 19012 9338 19068
rect 9338 19012 9394 19068
rect 9394 19012 9398 19068
rect 9334 19008 9398 19012
rect 14522 19068 14586 19072
rect 14522 19012 14526 19068
rect 14526 19012 14582 19068
rect 14582 19012 14586 19068
rect 14522 19008 14586 19012
rect 14602 19068 14666 19072
rect 14602 19012 14606 19068
rect 14606 19012 14662 19068
rect 14662 19012 14666 19068
rect 14602 19008 14666 19012
rect 14682 19068 14746 19072
rect 14682 19012 14686 19068
rect 14686 19012 14742 19068
rect 14742 19012 14746 19068
rect 14682 19008 14746 19012
rect 14762 19068 14826 19072
rect 14762 19012 14766 19068
rect 14766 19012 14822 19068
rect 14822 19012 14826 19068
rect 14762 19008 14826 19012
rect 19950 19068 20014 19072
rect 19950 19012 19954 19068
rect 19954 19012 20010 19068
rect 20010 19012 20014 19068
rect 19950 19008 20014 19012
rect 20030 19068 20094 19072
rect 20030 19012 20034 19068
rect 20034 19012 20090 19068
rect 20090 19012 20094 19068
rect 20030 19008 20094 19012
rect 20110 19068 20174 19072
rect 20110 19012 20114 19068
rect 20114 19012 20170 19068
rect 20170 19012 20174 19068
rect 20110 19008 20174 19012
rect 20190 19068 20254 19072
rect 20190 19012 20194 19068
rect 20194 19012 20250 19068
rect 20250 19012 20254 19068
rect 20190 19008 20254 19012
rect 6380 18524 6444 18528
rect 6380 18468 6384 18524
rect 6384 18468 6440 18524
rect 6440 18468 6444 18524
rect 6380 18464 6444 18468
rect 6460 18524 6524 18528
rect 6460 18468 6464 18524
rect 6464 18468 6520 18524
rect 6520 18468 6524 18524
rect 6460 18464 6524 18468
rect 6540 18524 6604 18528
rect 6540 18468 6544 18524
rect 6544 18468 6600 18524
rect 6600 18468 6604 18524
rect 6540 18464 6604 18468
rect 6620 18524 6684 18528
rect 6620 18468 6624 18524
rect 6624 18468 6680 18524
rect 6680 18468 6684 18524
rect 6620 18464 6684 18468
rect 11808 18524 11872 18528
rect 11808 18468 11812 18524
rect 11812 18468 11868 18524
rect 11868 18468 11872 18524
rect 11808 18464 11872 18468
rect 11888 18524 11952 18528
rect 11888 18468 11892 18524
rect 11892 18468 11948 18524
rect 11948 18468 11952 18524
rect 11888 18464 11952 18468
rect 11968 18524 12032 18528
rect 11968 18468 11972 18524
rect 11972 18468 12028 18524
rect 12028 18468 12032 18524
rect 11968 18464 12032 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 17316 18524 17380 18528
rect 17316 18468 17320 18524
rect 17320 18468 17376 18524
rect 17376 18468 17380 18524
rect 17316 18464 17380 18468
rect 17396 18524 17460 18528
rect 17396 18468 17400 18524
rect 17400 18468 17456 18524
rect 17456 18468 17460 18524
rect 17396 18464 17460 18468
rect 17476 18524 17540 18528
rect 17476 18468 17480 18524
rect 17480 18468 17536 18524
rect 17536 18468 17540 18524
rect 17476 18464 17540 18468
rect 22664 18524 22728 18528
rect 22664 18468 22668 18524
rect 22668 18468 22724 18524
rect 22724 18468 22728 18524
rect 22664 18464 22728 18468
rect 22744 18524 22808 18528
rect 22744 18468 22748 18524
rect 22748 18468 22804 18524
rect 22804 18468 22808 18524
rect 22744 18464 22808 18468
rect 22824 18524 22888 18528
rect 22824 18468 22828 18524
rect 22828 18468 22884 18524
rect 22884 18468 22888 18524
rect 22824 18464 22888 18468
rect 22904 18524 22968 18528
rect 22904 18468 22908 18524
rect 22908 18468 22964 18524
rect 22964 18468 22968 18524
rect 22904 18464 22968 18468
rect 3666 17980 3730 17984
rect 3666 17924 3670 17980
rect 3670 17924 3726 17980
rect 3726 17924 3730 17980
rect 3666 17920 3730 17924
rect 3746 17980 3810 17984
rect 3746 17924 3750 17980
rect 3750 17924 3806 17980
rect 3806 17924 3810 17980
rect 3746 17920 3810 17924
rect 3826 17980 3890 17984
rect 3826 17924 3830 17980
rect 3830 17924 3886 17980
rect 3886 17924 3890 17980
rect 3826 17920 3890 17924
rect 3906 17980 3970 17984
rect 3906 17924 3910 17980
rect 3910 17924 3966 17980
rect 3966 17924 3970 17980
rect 3906 17920 3970 17924
rect 9094 17980 9158 17984
rect 9094 17924 9098 17980
rect 9098 17924 9154 17980
rect 9154 17924 9158 17980
rect 9094 17920 9158 17924
rect 9174 17980 9238 17984
rect 9174 17924 9178 17980
rect 9178 17924 9234 17980
rect 9234 17924 9238 17980
rect 9174 17920 9238 17924
rect 9254 17980 9318 17984
rect 9254 17924 9258 17980
rect 9258 17924 9314 17980
rect 9314 17924 9318 17980
rect 9254 17920 9318 17924
rect 9334 17980 9398 17984
rect 9334 17924 9338 17980
rect 9338 17924 9394 17980
rect 9394 17924 9398 17980
rect 9334 17920 9398 17924
rect 14522 17980 14586 17984
rect 14522 17924 14526 17980
rect 14526 17924 14582 17980
rect 14582 17924 14586 17980
rect 14522 17920 14586 17924
rect 14602 17980 14666 17984
rect 14602 17924 14606 17980
rect 14606 17924 14662 17980
rect 14662 17924 14666 17980
rect 14602 17920 14666 17924
rect 14682 17980 14746 17984
rect 14682 17924 14686 17980
rect 14686 17924 14742 17980
rect 14742 17924 14746 17980
rect 14682 17920 14746 17924
rect 14762 17980 14826 17984
rect 14762 17924 14766 17980
rect 14766 17924 14822 17980
rect 14822 17924 14826 17980
rect 14762 17920 14826 17924
rect 19950 17980 20014 17984
rect 19950 17924 19954 17980
rect 19954 17924 20010 17980
rect 20010 17924 20014 17980
rect 19950 17920 20014 17924
rect 20030 17980 20094 17984
rect 20030 17924 20034 17980
rect 20034 17924 20090 17980
rect 20090 17924 20094 17980
rect 20030 17920 20094 17924
rect 20110 17980 20174 17984
rect 20110 17924 20114 17980
rect 20114 17924 20170 17980
rect 20170 17924 20174 17980
rect 20110 17920 20174 17924
rect 20190 17980 20254 17984
rect 20190 17924 20194 17980
rect 20194 17924 20250 17980
rect 20250 17924 20254 17980
rect 20190 17920 20254 17924
rect 6380 17436 6444 17440
rect 6380 17380 6384 17436
rect 6384 17380 6440 17436
rect 6440 17380 6444 17436
rect 6380 17376 6444 17380
rect 6460 17436 6524 17440
rect 6460 17380 6464 17436
rect 6464 17380 6520 17436
rect 6520 17380 6524 17436
rect 6460 17376 6524 17380
rect 6540 17436 6604 17440
rect 6540 17380 6544 17436
rect 6544 17380 6600 17436
rect 6600 17380 6604 17436
rect 6540 17376 6604 17380
rect 6620 17436 6684 17440
rect 6620 17380 6624 17436
rect 6624 17380 6680 17436
rect 6680 17380 6684 17436
rect 6620 17376 6684 17380
rect 11808 17436 11872 17440
rect 11808 17380 11812 17436
rect 11812 17380 11868 17436
rect 11868 17380 11872 17436
rect 11808 17376 11872 17380
rect 11888 17436 11952 17440
rect 11888 17380 11892 17436
rect 11892 17380 11948 17436
rect 11948 17380 11952 17436
rect 11888 17376 11952 17380
rect 11968 17436 12032 17440
rect 11968 17380 11972 17436
rect 11972 17380 12028 17436
rect 12028 17380 12032 17436
rect 11968 17376 12032 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 17316 17436 17380 17440
rect 17316 17380 17320 17436
rect 17320 17380 17376 17436
rect 17376 17380 17380 17436
rect 17316 17376 17380 17380
rect 17396 17436 17460 17440
rect 17396 17380 17400 17436
rect 17400 17380 17456 17436
rect 17456 17380 17460 17436
rect 17396 17376 17460 17380
rect 17476 17436 17540 17440
rect 17476 17380 17480 17436
rect 17480 17380 17536 17436
rect 17536 17380 17540 17436
rect 17476 17376 17540 17380
rect 22664 17436 22728 17440
rect 22664 17380 22668 17436
rect 22668 17380 22724 17436
rect 22724 17380 22728 17436
rect 22664 17376 22728 17380
rect 22744 17436 22808 17440
rect 22744 17380 22748 17436
rect 22748 17380 22804 17436
rect 22804 17380 22808 17436
rect 22744 17376 22808 17380
rect 22824 17436 22888 17440
rect 22824 17380 22828 17436
rect 22828 17380 22884 17436
rect 22884 17380 22888 17436
rect 22824 17376 22888 17380
rect 22904 17436 22968 17440
rect 22904 17380 22908 17436
rect 22908 17380 22964 17436
rect 22964 17380 22968 17436
rect 22904 17376 22968 17380
rect 3666 16892 3730 16896
rect 3666 16836 3670 16892
rect 3670 16836 3726 16892
rect 3726 16836 3730 16892
rect 3666 16832 3730 16836
rect 3746 16892 3810 16896
rect 3746 16836 3750 16892
rect 3750 16836 3806 16892
rect 3806 16836 3810 16892
rect 3746 16832 3810 16836
rect 3826 16892 3890 16896
rect 3826 16836 3830 16892
rect 3830 16836 3886 16892
rect 3886 16836 3890 16892
rect 3826 16832 3890 16836
rect 3906 16892 3970 16896
rect 3906 16836 3910 16892
rect 3910 16836 3966 16892
rect 3966 16836 3970 16892
rect 3906 16832 3970 16836
rect 9094 16892 9158 16896
rect 9094 16836 9098 16892
rect 9098 16836 9154 16892
rect 9154 16836 9158 16892
rect 9094 16832 9158 16836
rect 9174 16892 9238 16896
rect 9174 16836 9178 16892
rect 9178 16836 9234 16892
rect 9234 16836 9238 16892
rect 9174 16832 9238 16836
rect 9254 16892 9318 16896
rect 9254 16836 9258 16892
rect 9258 16836 9314 16892
rect 9314 16836 9318 16892
rect 9254 16832 9318 16836
rect 9334 16892 9398 16896
rect 9334 16836 9338 16892
rect 9338 16836 9394 16892
rect 9394 16836 9398 16892
rect 9334 16832 9398 16836
rect 14522 16892 14586 16896
rect 14522 16836 14526 16892
rect 14526 16836 14582 16892
rect 14582 16836 14586 16892
rect 14522 16832 14586 16836
rect 14602 16892 14666 16896
rect 14602 16836 14606 16892
rect 14606 16836 14662 16892
rect 14662 16836 14666 16892
rect 14602 16832 14666 16836
rect 14682 16892 14746 16896
rect 14682 16836 14686 16892
rect 14686 16836 14742 16892
rect 14742 16836 14746 16892
rect 14682 16832 14746 16836
rect 14762 16892 14826 16896
rect 14762 16836 14766 16892
rect 14766 16836 14822 16892
rect 14822 16836 14826 16892
rect 14762 16832 14826 16836
rect 19950 16892 20014 16896
rect 19950 16836 19954 16892
rect 19954 16836 20010 16892
rect 20010 16836 20014 16892
rect 19950 16832 20014 16836
rect 20030 16892 20094 16896
rect 20030 16836 20034 16892
rect 20034 16836 20090 16892
rect 20090 16836 20094 16892
rect 20030 16832 20094 16836
rect 20110 16892 20174 16896
rect 20110 16836 20114 16892
rect 20114 16836 20170 16892
rect 20170 16836 20174 16892
rect 20110 16832 20174 16836
rect 20190 16892 20254 16896
rect 20190 16836 20194 16892
rect 20194 16836 20250 16892
rect 20250 16836 20254 16892
rect 20190 16832 20254 16836
rect 6380 16348 6444 16352
rect 6380 16292 6384 16348
rect 6384 16292 6440 16348
rect 6440 16292 6444 16348
rect 6380 16288 6444 16292
rect 6460 16348 6524 16352
rect 6460 16292 6464 16348
rect 6464 16292 6520 16348
rect 6520 16292 6524 16348
rect 6460 16288 6524 16292
rect 6540 16348 6604 16352
rect 6540 16292 6544 16348
rect 6544 16292 6600 16348
rect 6600 16292 6604 16348
rect 6540 16288 6604 16292
rect 6620 16348 6684 16352
rect 6620 16292 6624 16348
rect 6624 16292 6680 16348
rect 6680 16292 6684 16348
rect 6620 16288 6684 16292
rect 11808 16348 11872 16352
rect 11808 16292 11812 16348
rect 11812 16292 11868 16348
rect 11868 16292 11872 16348
rect 11808 16288 11872 16292
rect 11888 16348 11952 16352
rect 11888 16292 11892 16348
rect 11892 16292 11948 16348
rect 11948 16292 11952 16348
rect 11888 16288 11952 16292
rect 11968 16348 12032 16352
rect 11968 16292 11972 16348
rect 11972 16292 12028 16348
rect 12028 16292 12032 16348
rect 11968 16288 12032 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 17316 16348 17380 16352
rect 17316 16292 17320 16348
rect 17320 16292 17376 16348
rect 17376 16292 17380 16348
rect 17316 16288 17380 16292
rect 17396 16348 17460 16352
rect 17396 16292 17400 16348
rect 17400 16292 17456 16348
rect 17456 16292 17460 16348
rect 17396 16288 17460 16292
rect 17476 16348 17540 16352
rect 17476 16292 17480 16348
rect 17480 16292 17536 16348
rect 17536 16292 17540 16348
rect 17476 16288 17540 16292
rect 22664 16348 22728 16352
rect 22664 16292 22668 16348
rect 22668 16292 22724 16348
rect 22724 16292 22728 16348
rect 22664 16288 22728 16292
rect 22744 16348 22808 16352
rect 22744 16292 22748 16348
rect 22748 16292 22804 16348
rect 22804 16292 22808 16348
rect 22744 16288 22808 16292
rect 22824 16348 22888 16352
rect 22824 16292 22828 16348
rect 22828 16292 22884 16348
rect 22884 16292 22888 16348
rect 22824 16288 22888 16292
rect 22904 16348 22968 16352
rect 22904 16292 22908 16348
rect 22908 16292 22964 16348
rect 22964 16292 22968 16348
rect 22904 16288 22968 16292
rect 3666 15804 3730 15808
rect 3666 15748 3670 15804
rect 3670 15748 3726 15804
rect 3726 15748 3730 15804
rect 3666 15744 3730 15748
rect 3746 15804 3810 15808
rect 3746 15748 3750 15804
rect 3750 15748 3806 15804
rect 3806 15748 3810 15804
rect 3746 15744 3810 15748
rect 3826 15804 3890 15808
rect 3826 15748 3830 15804
rect 3830 15748 3886 15804
rect 3886 15748 3890 15804
rect 3826 15744 3890 15748
rect 3906 15804 3970 15808
rect 3906 15748 3910 15804
rect 3910 15748 3966 15804
rect 3966 15748 3970 15804
rect 3906 15744 3970 15748
rect 9094 15804 9158 15808
rect 9094 15748 9098 15804
rect 9098 15748 9154 15804
rect 9154 15748 9158 15804
rect 9094 15744 9158 15748
rect 9174 15804 9238 15808
rect 9174 15748 9178 15804
rect 9178 15748 9234 15804
rect 9234 15748 9238 15804
rect 9174 15744 9238 15748
rect 9254 15804 9318 15808
rect 9254 15748 9258 15804
rect 9258 15748 9314 15804
rect 9314 15748 9318 15804
rect 9254 15744 9318 15748
rect 9334 15804 9398 15808
rect 9334 15748 9338 15804
rect 9338 15748 9394 15804
rect 9394 15748 9398 15804
rect 9334 15744 9398 15748
rect 14522 15804 14586 15808
rect 14522 15748 14526 15804
rect 14526 15748 14582 15804
rect 14582 15748 14586 15804
rect 14522 15744 14586 15748
rect 14602 15804 14666 15808
rect 14602 15748 14606 15804
rect 14606 15748 14662 15804
rect 14662 15748 14666 15804
rect 14602 15744 14666 15748
rect 14682 15804 14746 15808
rect 14682 15748 14686 15804
rect 14686 15748 14742 15804
rect 14742 15748 14746 15804
rect 14682 15744 14746 15748
rect 14762 15804 14826 15808
rect 14762 15748 14766 15804
rect 14766 15748 14822 15804
rect 14822 15748 14826 15804
rect 14762 15744 14826 15748
rect 19950 15804 20014 15808
rect 19950 15748 19954 15804
rect 19954 15748 20010 15804
rect 20010 15748 20014 15804
rect 19950 15744 20014 15748
rect 20030 15804 20094 15808
rect 20030 15748 20034 15804
rect 20034 15748 20090 15804
rect 20090 15748 20094 15804
rect 20030 15744 20094 15748
rect 20110 15804 20174 15808
rect 20110 15748 20114 15804
rect 20114 15748 20170 15804
rect 20170 15748 20174 15804
rect 20110 15744 20174 15748
rect 20190 15804 20254 15808
rect 20190 15748 20194 15804
rect 20194 15748 20250 15804
rect 20250 15748 20254 15804
rect 20190 15744 20254 15748
rect 6380 15260 6444 15264
rect 6380 15204 6384 15260
rect 6384 15204 6440 15260
rect 6440 15204 6444 15260
rect 6380 15200 6444 15204
rect 6460 15260 6524 15264
rect 6460 15204 6464 15260
rect 6464 15204 6520 15260
rect 6520 15204 6524 15260
rect 6460 15200 6524 15204
rect 6540 15260 6604 15264
rect 6540 15204 6544 15260
rect 6544 15204 6600 15260
rect 6600 15204 6604 15260
rect 6540 15200 6604 15204
rect 6620 15260 6684 15264
rect 6620 15204 6624 15260
rect 6624 15204 6680 15260
rect 6680 15204 6684 15260
rect 6620 15200 6684 15204
rect 11808 15260 11872 15264
rect 11808 15204 11812 15260
rect 11812 15204 11868 15260
rect 11868 15204 11872 15260
rect 11808 15200 11872 15204
rect 11888 15260 11952 15264
rect 11888 15204 11892 15260
rect 11892 15204 11948 15260
rect 11948 15204 11952 15260
rect 11888 15200 11952 15204
rect 11968 15260 12032 15264
rect 11968 15204 11972 15260
rect 11972 15204 12028 15260
rect 12028 15204 12032 15260
rect 11968 15200 12032 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 17316 15260 17380 15264
rect 17316 15204 17320 15260
rect 17320 15204 17376 15260
rect 17376 15204 17380 15260
rect 17316 15200 17380 15204
rect 17396 15260 17460 15264
rect 17396 15204 17400 15260
rect 17400 15204 17456 15260
rect 17456 15204 17460 15260
rect 17396 15200 17460 15204
rect 17476 15260 17540 15264
rect 17476 15204 17480 15260
rect 17480 15204 17536 15260
rect 17536 15204 17540 15260
rect 17476 15200 17540 15204
rect 22664 15260 22728 15264
rect 22664 15204 22668 15260
rect 22668 15204 22724 15260
rect 22724 15204 22728 15260
rect 22664 15200 22728 15204
rect 22744 15260 22808 15264
rect 22744 15204 22748 15260
rect 22748 15204 22804 15260
rect 22804 15204 22808 15260
rect 22744 15200 22808 15204
rect 22824 15260 22888 15264
rect 22824 15204 22828 15260
rect 22828 15204 22884 15260
rect 22884 15204 22888 15260
rect 22824 15200 22888 15204
rect 22904 15260 22968 15264
rect 22904 15204 22908 15260
rect 22908 15204 22964 15260
rect 22964 15204 22968 15260
rect 22904 15200 22968 15204
rect 3666 14716 3730 14720
rect 3666 14660 3670 14716
rect 3670 14660 3726 14716
rect 3726 14660 3730 14716
rect 3666 14656 3730 14660
rect 3746 14716 3810 14720
rect 3746 14660 3750 14716
rect 3750 14660 3806 14716
rect 3806 14660 3810 14716
rect 3746 14656 3810 14660
rect 3826 14716 3890 14720
rect 3826 14660 3830 14716
rect 3830 14660 3886 14716
rect 3886 14660 3890 14716
rect 3826 14656 3890 14660
rect 3906 14716 3970 14720
rect 3906 14660 3910 14716
rect 3910 14660 3966 14716
rect 3966 14660 3970 14716
rect 3906 14656 3970 14660
rect 9094 14716 9158 14720
rect 9094 14660 9098 14716
rect 9098 14660 9154 14716
rect 9154 14660 9158 14716
rect 9094 14656 9158 14660
rect 9174 14716 9238 14720
rect 9174 14660 9178 14716
rect 9178 14660 9234 14716
rect 9234 14660 9238 14716
rect 9174 14656 9238 14660
rect 9254 14716 9318 14720
rect 9254 14660 9258 14716
rect 9258 14660 9314 14716
rect 9314 14660 9318 14716
rect 9254 14656 9318 14660
rect 9334 14716 9398 14720
rect 9334 14660 9338 14716
rect 9338 14660 9394 14716
rect 9394 14660 9398 14716
rect 9334 14656 9398 14660
rect 14522 14716 14586 14720
rect 14522 14660 14526 14716
rect 14526 14660 14582 14716
rect 14582 14660 14586 14716
rect 14522 14656 14586 14660
rect 14602 14716 14666 14720
rect 14602 14660 14606 14716
rect 14606 14660 14662 14716
rect 14662 14660 14666 14716
rect 14602 14656 14666 14660
rect 14682 14716 14746 14720
rect 14682 14660 14686 14716
rect 14686 14660 14742 14716
rect 14742 14660 14746 14716
rect 14682 14656 14746 14660
rect 14762 14716 14826 14720
rect 14762 14660 14766 14716
rect 14766 14660 14822 14716
rect 14822 14660 14826 14716
rect 14762 14656 14826 14660
rect 19950 14716 20014 14720
rect 19950 14660 19954 14716
rect 19954 14660 20010 14716
rect 20010 14660 20014 14716
rect 19950 14656 20014 14660
rect 20030 14716 20094 14720
rect 20030 14660 20034 14716
rect 20034 14660 20090 14716
rect 20090 14660 20094 14716
rect 20030 14656 20094 14660
rect 20110 14716 20174 14720
rect 20110 14660 20114 14716
rect 20114 14660 20170 14716
rect 20170 14660 20174 14716
rect 20110 14656 20174 14660
rect 20190 14716 20254 14720
rect 20190 14660 20194 14716
rect 20194 14660 20250 14716
rect 20250 14660 20254 14716
rect 20190 14656 20254 14660
rect 6380 14172 6444 14176
rect 6380 14116 6384 14172
rect 6384 14116 6440 14172
rect 6440 14116 6444 14172
rect 6380 14112 6444 14116
rect 6460 14172 6524 14176
rect 6460 14116 6464 14172
rect 6464 14116 6520 14172
rect 6520 14116 6524 14172
rect 6460 14112 6524 14116
rect 6540 14172 6604 14176
rect 6540 14116 6544 14172
rect 6544 14116 6600 14172
rect 6600 14116 6604 14172
rect 6540 14112 6604 14116
rect 6620 14172 6684 14176
rect 6620 14116 6624 14172
rect 6624 14116 6680 14172
rect 6680 14116 6684 14172
rect 6620 14112 6684 14116
rect 11808 14172 11872 14176
rect 11808 14116 11812 14172
rect 11812 14116 11868 14172
rect 11868 14116 11872 14172
rect 11808 14112 11872 14116
rect 11888 14172 11952 14176
rect 11888 14116 11892 14172
rect 11892 14116 11948 14172
rect 11948 14116 11952 14172
rect 11888 14112 11952 14116
rect 11968 14172 12032 14176
rect 11968 14116 11972 14172
rect 11972 14116 12028 14172
rect 12028 14116 12032 14172
rect 11968 14112 12032 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 17316 14172 17380 14176
rect 17316 14116 17320 14172
rect 17320 14116 17376 14172
rect 17376 14116 17380 14172
rect 17316 14112 17380 14116
rect 17396 14172 17460 14176
rect 17396 14116 17400 14172
rect 17400 14116 17456 14172
rect 17456 14116 17460 14172
rect 17396 14112 17460 14116
rect 17476 14172 17540 14176
rect 17476 14116 17480 14172
rect 17480 14116 17536 14172
rect 17536 14116 17540 14172
rect 17476 14112 17540 14116
rect 22664 14172 22728 14176
rect 22664 14116 22668 14172
rect 22668 14116 22724 14172
rect 22724 14116 22728 14172
rect 22664 14112 22728 14116
rect 22744 14172 22808 14176
rect 22744 14116 22748 14172
rect 22748 14116 22804 14172
rect 22804 14116 22808 14172
rect 22744 14112 22808 14116
rect 22824 14172 22888 14176
rect 22824 14116 22828 14172
rect 22828 14116 22884 14172
rect 22884 14116 22888 14172
rect 22824 14112 22888 14116
rect 22904 14172 22968 14176
rect 22904 14116 22908 14172
rect 22908 14116 22964 14172
rect 22964 14116 22968 14172
rect 22904 14112 22968 14116
rect 3666 13628 3730 13632
rect 3666 13572 3670 13628
rect 3670 13572 3726 13628
rect 3726 13572 3730 13628
rect 3666 13568 3730 13572
rect 3746 13628 3810 13632
rect 3746 13572 3750 13628
rect 3750 13572 3806 13628
rect 3806 13572 3810 13628
rect 3746 13568 3810 13572
rect 3826 13628 3890 13632
rect 3826 13572 3830 13628
rect 3830 13572 3886 13628
rect 3886 13572 3890 13628
rect 3826 13568 3890 13572
rect 3906 13628 3970 13632
rect 3906 13572 3910 13628
rect 3910 13572 3966 13628
rect 3966 13572 3970 13628
rect 3906 13568 3970 13572
rect 9094 13628 9158 13632
rect 9094 13572 9098 13628
rect 9098 13572 9154 13628
rect 9154 13572 9158 13628
rect 9094 13568 9158 13572
rect 9174 13628 9238 13632
rect 9174 13572 9178 13628
rect 9178 13572 9234 13628
rect 9234 13572 9238 13628
rect 9174 13568 9238 13572
rect 9254 13628 9318 13632
rect 9254 13572 9258 13628
rect 9258 13572 9314 13628
rect 9314 13572 9318 13628
rect 9254 13568 9318 13572
rect 9334 13628 9398 13632
rect 9334 13572 9338 13628
rect 9338 13572 9394 13628
rect 9394 13572 9398 13628
rect 9334 13568 9398 13572
rect 14522 13628 14586 13632
rect 14522 13572 14526 13628
rect 14526 13572 14582 13628
rect 14582 13572 14586 13628
rect 14522 13568 14586 13572
rect 14602 13628 14666 13632
rect 14602 13572 14606 13628
rect 14606 13572 14662 13628
rect 14662 13572 14666 13628
rect 14602 13568 14666 13572
rect 14682 13628 14746 13632
rect 14682 13572 14686 13628
rect 14686 13572 14742 13628
rect 14742 13572 14746 13628
rect 14682 13568 14746 13572
rect 14762 13628 14826 13632
rect 14762 13572 14766 13628
rect 14766 13572 14822 13628
rect 14822 13572 14826 13628
rect 14762 13568 14826 13572
rect 19950 13628 20014 13632
rect 19950 13572 19954 13628
rect 19954 13572 20010 13628
rect 20010 13572 20014 13628
rect 19950 13568 20014 13572
rect 20030 13628 20094 13632
rect 20030 13572 20034 13628
rect 20034 13572 20090 13628
rect 20090 13572 20094 13628
rect 20030 13568 20094 13572
rect 20110 13628 20174 13632
rect 20110 13572 20114 13628
rect 20114 13572 20170 13628
rect 20170 13572 20174 13628
rect 20110 13568 20174 13572
rect 20190 13628 20254 13632
rect 20190 13572 20194 13628
rect 20194 13572 20250 13628
rect 20250 13572 20254 13628
rect 20190 13568 20254 13572
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 11808 13084 11872 13088
rect 11808 13028 11812 13084
rect 11812 13028 11868 13084
rect 11868 13028 11872 13084
rect 11808 13024 11872 13028
rect 11888 13084 11952 13088
rect 11888 13028 11892 13084
rect 11892 13028 11948 13084
rect 11948 13028 11952 13084
rect 11888 13024 11952 13028
rect 11968 13084 12032 13088
rect 11968 13028 11972 13084
rect 11972 13028 12028 13084
rect 12028 13028 12032 13084
rect 11968 13024 12032 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 17316 13084 17380 13088
rect 17316 13028 17320 13084
rect 17320 13028 17376 13084
rect 17376 13028 17380 13084
rect 17316 13024 17380 13028
rect 17396 13084 17460 13088
rect 17396 13028 17400 13084
rect 17400 13028 17456 13084
rect 17456 13028 17460 13084
rect 17396 13024 17460 13028
rect 17476 13084 17540 13088
rect 17476 13028 17480 13084
rect 17480 13028 17536 13084
rect 17536 13028 17540 13084
rect 17476 13024 17540 13028
rect 22664 13084 22728 13088
rect 22664 13028 22668 13084
rect 22668 13028 22724 13084
rect 22724 13028 22728 13084
rect 22664 13024 22728 13028
rect 22744 13084 22808 13088
rect 22744 13028 22748 13084
rect 22748 13028 22804 13084
rect 22804 13028 22808 13084
rect 22744 13024 22808 13028
rect 22824 13084 22888 13088
rect 22824 13028 22828 13084
rect 22828 13028 22884 13084
rect 22884 13028 22888 13084
rect 22824 13024 22888 13028
rect 22904 13084 22968 13088
rect 22904 13028 22908 13084
rect 22908 13028 22964 13084
rect 22964 13028 22968 13084
rect 22904 13024 22968 13028
rect 3666 12540 3730 12544
rect 3666 12484 3670 12540
rect 3670 12484 3726 12540
rect 3726 12484 3730 12540
rect 3666 12480 3730 12484
rect 3746 12540 3810 12544
rect 3746 12484 3750 12540
rect 3750 12484 3806 12540
rect 3806 12484 3810 12540
rect 3746 12480 3810 12484
rect 3826 12540 3890 12544
rect 3826 12484 3830 12540
rect 3830 12484 3886 12540
rect 3886 12484 3890 12540
rect 3826 12480 3890 12484
rect 3906 12540 3970 12544
rect 3906 12484 3910 12540
rect 3910 12484 3966 12540
rect 3966 12484 3970 12540
rect 3906 12480 3970 12484
rect 9094 12540 9158 12544
rect 9094 12484 9098 12540
rect 9098 12484 9154 12540
rect 9154 12484 9158 12540
rect 9094 12480 9158 12484
rect 9174 12540 9238 12544
rect 9174 12484 9178 12540
rect 9178 12484 9234 12540
rect 9234 12484 9238 12540
rect 9174 12480 9238 12484
rect 9254 12540 9318 12544
rect 9254 12484 9258 12540
rect 9258 12484 9314 12540
rect 9314 12484 9318 12540
rect 9254 12480 9318 12484
rect 9334 12540 9398 12544
rect 9334 12484 9338 12540
rect 9338 12484 9394 12540
rect 9394 12484 9398 12540
rect 9334 12480 9398 12484
rect 14522 12540 14586 12544
rect 14522 12484 14526 12540
rect 14526 12484 14582 12540
rect 14582 12484 14586 12540
rect 14522 12480 14586 12484
rect 14602 12540 14666 12544
rect 14602 12484 14606 12540
rect 14606 12484 14662 12540
rect 14662 12484 14666 12540
rect 14602 12480 14666 12484
rect 14682 12540 14746 12544
rect 14682 12484 14686 12540
rect 14686 12484 14742 12540
rect 14742 12484 14746 12540
rect 14682 12480 14746 12484
rect 14762 12540 14826 12544
rect 14762 12484 14766 12540
rect 14766 12484 14822 12540
rect 14822 12484 14826 12540
rect 14762 12480 14826 12484
rect 19950 12540 20014 12544
rect 19950 12484 19954 12540
rect 19954 12484 20010 12540
rect 20010 12484 20014 12540
rect 19950 12480 20014 12484
rect 20030 12540 20094 12544
rect 20030 12484 20034 12540
rect 20034 12484 20090 12540
rect 20090 12484 20094 12540
rect 20030 12480 20094 12484
rect 20110 12540 20174 12544
rect 20110 12484 20114 12540
rect 20114 12484 20170 12540
rect 20170 12484 20174 12540
rect 20110 12480 20174 12484
rect 20190 12540 20254 12544
rect 20190 12484 20194 12540
rect 20194 12484 20250 12540
rect 20250 12484 20254 12540
rect 20190 12480 20254 12484
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 11808 11996 11872 12000
rect 11808 11940 11812 11996
rect 11812 11940 11868 11996
rect 11868 11940 11872 11996
rect 11808 11936 11872 11940
rect 11888 11996 11952 12000
rect 11888 11940 11892 11996
rect 11892 11940 11948 11996
rect 11948 11940 11952 11996
rect 11888 11936 11952 11940
rect 11968 11996 12032 12000
rect 11968 11940 11972 11996
rect 11972 11940 12028 11996
rect 12028 11940 12032 11996
rect 11968 11936 12032 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 17316 11996 17380 12000
rect 17316 11940 17320 11996
rect 17320 11940 17376 11996
rect 17376 11940 17380 11996
rect 17316 11936 17380 11940
rect 17396 11996 17460 12000
rect 17396 11940 17400 11996
rect 17400 11940 17456 11996
rect 17456 11940 17460 11996
rect 17396 11936 17460 11940
rect 17476 11996 17540 12000
rect 17476 11940 17480 11996
rect 17480 11940 17536 11996
rect 17536 11940 17540 11996
rect 17476 11936 17540 11940
rect 22664 11996 22728 12000
rect 22664 11940 22668 11996
rect 22668 11940 22724 11996
rect 22724 11940 22728 11996
rect 22664 11936 22728 11940
rect 22744 11996 22808 12000
rect 22744 11940 22748 11996
rect 22748 11940 22804 11996
rect 22804 11940 22808 11996
rect 22744 11936 22808 11940
rect 22824 11996 22888 12000
rect 22824 11940 22828 11996
rect 22828 11940 22884 11996
rect 22884 11940 22888 11996
rect 22824 11936 22888 11940
rect 22904 11996 22968 12000
rect 22904 11940 22908 11996
rect 22908 11940 22964 11996
rect 22964 11940 22968 11996
rect 22904 11936 22968 11940
rect 3666 11452 3730 11456
rect 3666 11396 3670 11452
rect 3670 11396 3726 11452
rect 3726 11396 3730 11452
rect 3666 11392 3730 11396
rect 3746 11452 3810 11456
rect 3746 11396 3750 11452
rect 3750 11396 3806 11452
rect 3806 11396 3810 11452
rect 3746 11392 3810 11396
rect 3826 11452 3890 11456
rect 3826 11396 3830 11452
rect 3830 11396 3886 11452
rect 3886 11396 3890 11452
rect 3826 11392 3890 11396
rect 3906 11452 3970 11456
rect 3906 11396 3910 11452
rect 3910 11396 3966 11452
rect 3966 11396 3970 11452
rect 3906 11392 3970 11396
rect 9094 11452 9158 11456
rect 9094 11396 9098 11452
rect 9098 11396 9154 11452
rect 9154 11396 9158 11452
rect 9094 11392 9158 11396
rect 9174 11452 9238 11456
rect 9174 11396 9178 11452
rect 9178 11396 9234 11452
rect 9234 11396 9238 11452
rect 9174 11392 9238 11396
rect 9254 11452 9318 11456
rect 9254 11396 9258 11452
rect 9258 11396 9314 11452
rect 9314 11396 9318 11452
rect 9254 11392 9318 11396
rect 9334 11452 9398 11456
rect 9334 11396 9338 11452
rect 9338 11396 9394 11452
rect 9394 11396 9398 11452
rect 9334 11392 9398 11396
rect 14522 11452 14586 11456
rect 14522 11396 14526 11452
rect 14526 11396 14582 11452
rect 14582 11396 14586 11452
rect 14522 11392 14586 11396
rect 14602 11452 14666 11456
rect 14602 11396 14606 11452
rect 14606 11396 14662 11452
rect 14662 11396 14666 11452
rect 14602 11392 14666 11396
rect 14682 11452 14746 11456
rect 14682 11396 14686 11452
rect 14686 11396 14742 11452
rect 14742 11396 14746 11452
rect 14682 11392 14746 11396
rect 14762 11452 14826 11456
rect 14762 11396 14766 11452
rect 14766 11396 14822 11452
rect 14822 11396 14826 11452
rect 14762 11392 14826 11396
rect 19950 11452 20014 11456
rect 19950 11396 19954 11452
rect 19954 11396 20010 11452
rect 20010 11396 20014 11452
rect 19950 11392 20014 11396
rect 20030 11452 20094 11456
rect 20030 11396 20034 11452
rect 20034 11396 20090 11452
rect 20090 11396 20094 11452
rect 20030 11392 20094 11396
rect 20110 11452 20174 11456
rect 20110 11396 20114 11452
rect 20114 11396 20170 11452
rect 20170 11396 20174 11452
rect 20110 11392 20174 11396
rect 20190 11452 20254 11456
rect 20190 11396 20194 11452
rect 20194 11396 20250 11452
rect 20250 11396 20254 11452
rect 20190 11392 20254 11396
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 11808 10908 11872 10912
rect 11808 10852 11812 10908
rect 11812 10852 11868 10908
rect 11868 10852 11872 10908
rect 11808 10848 11872 10852
rect 11888 10908 11952 10912
rect 11888 10852 11892 10908
rect 11892 10852 11948 10908
rect 11948 10852 11952 10908
rect 11888 10848 11952 10852
rect 11968 10908 12032 10912
rect 11968 10852 11972 10908
rect 11972 10852 12028 10908
rect 12028 10852 12032 10908
rect 11968 10848 12032 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 17316 10908 17380 10912
rect 17316 10852 17320 10908
rect 17320 10852 17376 10908
rect 17376 10852 17380 10908
rect 17316 10848 17380 10852
rect 17396 10908 17460 10912
rect 17396 10852 17400 10908
rect 17400 10852 17456 10908
rect 17456 10852 17460 10908
rect 17396 10848 17460 10852
rect 17476 10908 17540 10912
rect 17476 10852 17480 10908
rect 17480 10852 17536 10908
rect 17536 10852 17540 10908
rect 17476 10848 17540 10852
rect 22664 10908 22728 10912
rect 22664 10852 22668 10908
rect 22668 10852 22724 10908
rect 22724 10852 22728 10908
rect 22664 10848 22728 10852
rect 22744 10908 22808 10912
rect 22744 10852 22748 10908
rect 22748 10852 22804 10908
rect 22804 10852 22808 10908
rect 22744 10848 22808 10852
rect 22824 10908 22888 10912
rect 22824 10852 22828 10908
rect 22828 10852 22884 10908
rect 22884 10852 22888 10908
rect 22824 10848 22888 10852
rect 22904 10908 22968 10912
rect 22904 10852 22908 10908
rect 22908 10852 22964 10908
rect 22964 10852 22968 10908
rect 22904 10848 22968 10852
rect 3666 10364 3730 10368
rect 3666 10308 3670 10364
rect 3670 10308 3726 10364
rect 3726 10308 3730 10364
rect 3666 10304 3730 10308
rect 3746 10364 3810 10368
rect 3746 10308 3750 10364
rect 3750 10308 3806 10364
rect 3806 10308 3810 10364
rect 3746 10304 3810 10308
rect 3826 10364 3890 10368
rect 3826 10308 3830 10364
rect 3830 10308 3886 10364
rect 3886 10308 3890 10364
rect 3826 10304 3890 10308
rect 3906 10364 3970 10368
rect 3906 10308 3910 10364
rect 3910 10308 3966 10364
rect 3966 10308 3970 10364
rect 3906 10304 3970 10308
rect 9094 10364 9158 10368
rect 9094 10308 9098 10364
rect 9098 10308 9154 10364
rect 9154 10308 9158 10364
rect 9094 10304 9158 10308
rect 9174 10364 9238 10368
rect 9174 10308 9178 10364
rect 9178 10308 9234 10364
rect 9234 10308 9238 10364
rect 9174 10304 9238 10308
rect 9254 10364 9318 10368
rect 9254 10308 9258 10364
rect 9258 10308 9314 10364
rect 9314 10308 9318 10364
rect 9254 10304 9318 10308
rect 9334 10364 9398 10368
rect 9334 10308 9338 10364
rect 9338 10308 9394 10364
rect 9394 10308 9398 10364
rect 9334 10304 9398 10308
rect 14522 10364 14586 10368
rect 14522 10308 14526 10364
rect 14526 10308 14582 10364
rect 14582 10308 14586 10364
rect 14522 10304 14586 10308
rect 14602 10364 14666 10368
rect 14602 10308 14606 10364
rect 14606 10308 14662 10364
rect 14662 10308 14666 10364
rect 14602 10304 14666 10308
rect 14682 10364 14746 10368
rect 14682 10308 14686 10364
rect 14686 10308 14742 10364
rect 14742 10308 14746 10364
rect 14682 10304 14746 10308
rect 14762 10364 14826 10368
rect 14762 10308 14766 10364
rect 14766 10308 14822 10364
rect 14822 10308 14826 10364
rect 14762 10304 14826 10308
rect 19950 10364 20014 10368
rect 19950 10308 19954 10364
rect 19954 10308 20010 10364
rect 20010 10308 20014 10364
rect 19950 10304 20014 10308
rect 20030 10364 20094 10368
rect 20030 10308 20034 10364
rect 20034 10308 20090 10364
rect 20090 10308 20094 10364
rect 20030 10304 20094 10308
rect 20110 10364 20174 10368
rect 20110 10308 20114 10364
rect 20114 10308 20170 10364
rect 20170 10308 20174 10364
rect 20110 10304 20174 10308
rect 20190 10364 20254 10368
rect 20190 10308 20194 10364
rect 20194 10308 20250 10364
rect 20250 10308 20254 10364
rect 20190 10304 20254 10308
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 11808 9820 11872 9824
rect 11808 9764 11812 9820
rect 11812 9764 11868 9820
rect 11868 9764 11872 9820
rect 11808 9760 11872 9764
rect 11888 9820 11952 9824
rect 11888 9764 11892 9820
rect 11892 9764 11948 9820
rect 11948 9764 11952 9820
rect 11888 9760 11952 9764
rect 11968 9820 12032 9824
rect 11968 9764 11972 9820
rect 11972 9764 12028 9820
rect 12028 9764 12032 9820
rect 11968 9760 12032 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 17316 9820 17380 9824
rect 17316 9764 17320 9820
rect 17320 9764 17376 9820
rect 17376 9764 17380 9820
rect 17316 9760 17380 9764
rect 17396 9820 17460 9824
rect 17396 9764 17400 9820
rect 17400 9764 17456 9820
rect 17456 9764 17460 9820
rect 17396 9760 17460 9764
rect 17476 9820 17540 9824
rect 17476 9764 17480 9820
rect 17480 9764 17536 9820
rect 17536 9764 17540 9820
rect 17476 9760 17540 9764
rect 22664 9820 22728 9824
rect 22664 9764 22668 9820
rect 22668 9764 22724 9820
rect 22724 9764 22728 9820
rect 22664 9760 22728 9764
rect 22744 9820 22808 9824
rect 22744 9764 22748 9820
rect 22748 9764 22804 9820
rect 22804 9764 22808 9820
rect 22744 9760 22808 9764
rect 22824 9820 22888 9824
rect 22824 9764 22828 9820
rect 22828 9764 22884 9820
rect 22884 9764 22888 9820
rect 22824 9760 22888 9764
rect 22904 9820 22968 9824
rect 22904 9764 22908 9820
rect 22908 9764 22964 9820
rect 22964 9764 22968 9820
rect 22904 9760 22968 9764
rect 3666 9276 3730 9280
rect 3666 9220 3670 9276
rect 3670 9220 3726 9276
rect 3726 9220 3730 9276
rect 3666 9216 3730 9220
rect 3746 9276 3810 9280
rect 3746 9220 3750 9276
rect 3750 9220 3806 9276
rect 3806 9220 3810 9276
rect 3746 9216 3810 9220
rect 3826 9276 3890 9280
rect 3826 9220 3830 9276
rect 3830 9220 3886 9276
rect 3886 9220 3890 9276
rect 3826 9216 3890 9220
rect 3906 9276 3970 9280
rect 3906 9220 3910 9276
rect 3910 9220 3966 9276
rect 3966 9220 3970 9276
rect 3906 9216 3970 9220
rect 9094 9276 9158 9280
rect 9094 9220 9098 9276
rect 9098 9220 9154 9276
rect 9154 9220 9158 9276
rect 9094 9216 9158 9220
rect 9174 9276 9238 9280
rect 9174 9220 9178 9276
rect 9178 9220 9234 9276
rect 9234 9220 9238 9276
rect 9174 9216 9238 9220
rect 9254 9276 9318 9280
rect 9254 9220 9258 9276
rect 9258 9220 9314 9276
rect 9314 9220 9318 9276
rect 9254 9216 9318 9220
rect 9334 9276 9398 9280
rect 9334 9220 9338 9276
rect 9338 9220 9394 9276
rect 9394 9220 9398 9276
rect 9334 9216 9398 9220
rect 14522 9276 14586 9280
rect 14522 9220 14526 9276
rect 14526 9220 14582 9276
rect 14582 9220 14586 9276
rect 14522 9216 14586 9220
rect 14602 9276 14666 9280
rect 14602 9220 14606 9276
rect 14606 9220 14662 9276
rect 14662 9220 14666 9276
rect 14602 9216 14666 9220
rect 14682 9276 14746 9280
rect 14682 9220 14686 9276
rect 14686 9220 14742 9276
rect 14742 9220 14746 9276
rect 14682 9216 14746 9220
rect 14762 9276 14826 9280
rect 14762 9220 14766 9276
rect 14766 9220 14822 9276
rect 14822 9220 14826 9276
rect 14762 9216 14826 9220
rect 19950 9276 20014 9280
rect 19950 9220 19954 9276
rect 19954 9220 20010 9276
rect 20010 9220 20014 9276
rect 19950 9216 20014 9220
rect 20030 9276 20094 9280
rect 20030 9220 20034 9276
rect 20034 9220 20090 9276
rect 20090 9220 20094 9276
rect 20030 9216 20094 9220
rect 20110 9276 20174 9280
rect 20110 9220 20114 9276
rect 20114 9220 20170 9276
rect 20170 9220 20174 9276
rect 20110 9216 20174 9220
rect 20190 9276 20254 9280
rect 20190 9220 20194 9276
rect 20194 9220 20250 9276
rect 20250 9220 20254 9276
rect 20190 9216 20254 9220
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 11808 8732 11872 8736
rect 11808 8676 11812 8732
rect 11812 8676 11868 8732
rect 11868 8676 11872 8732
rect 11808 8672 11872 8676
rect 11888 8732 11952 8736
rect 11888 8676 11892 8732
rect 11892 8676 11948 8732
rect 11948 8676 11952 8732
rect 11888 8672 11952 8676
rect 11968 8732 12032 8736
rect 11968 8676 11972 8732
rect 11972 8676 12028 8732
rect 12028 8676 12032 8732
rect 11968 8672 12032 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 17316 8732 17380 8736
rect 17316 8676 17320 8732
rect 17320 8676 17376 8732
rect 17376 8676 17380 8732
rect 17316 8672 17380 8676
rect 17396 8732 17460 8736
rect 17396 8676 17400 8732
rect 17400 8676 17456 8732
rect 17456 8676 17460 8732
rect 17396 8672 17460 8676
rect 17476 8732 17540 8736
rect 17476 8676 17480 8732
rect 17480 8676 17536 8732
rect 17536 8676 17540 8732
rect 17476 8672 17540 8676
rect 22664 8732 22728 8736
rect 22664 8676 22668 8732
rect 22668 8676 22724 8732
rect 22724 8676 22728 8732
rect 22664 8672 22728 8676
rect 22744 8732 22808 8736
rect 22744 8676 22748 8732
rect 22748 8676 22804 8732
rect 22804 8676 22808 8732
rect 22744 8672 22808 8676
rect 22824 8732 22888 8736
rect 22824 8676 22828 8732
rect 22828 8676 22884 8732
rect 22884 8676 22888 8732
rect 22824 8672 22888 8676
rect 22904 8732 22968 8736
rect 22904 8676 22908 8732
rect 22908 8676 22964 8732
rect 22964 8676 22968 8732
rect 22904 8672 22968 8676
rect 3666 8188 3730 8192
rect 3666 8132 3670 8188
rect 3670 8132 3726 8188
rect 3726 8132 3730 8188
rect 3666 8128 3730 8132
rect 3746 8188 3810 8192
rect 3746 8132 3750 8188
rect 3750 8132 3806 8188
rect 3806 8132 3810 8188
rect 3746 8128 3810 8132
rect 3826 8188 3890 8192
rect 3826 8132 3830 8188
rect 3830 8132 3886 8188
rect 3886 8132 3890 8188
rect 3826 8128 3890 8132
rect 3906 8188 3970 8192
rect 3906 8132 3910 8188
rect 3910 8132 3966 8188
rect 3966 8132 3970 8188
rect 3906 8128 3970 8132
rect 9094 8188 9158 8192
rect 9094 8132 9098 8188
rect 9098 8132 9154 8188
rect 9154 8132 9158 8188
rect 9094 8128 9158 8132
rect 9174 8188 9238 8192
rect 9174 8132 9178 8188
rect 9178 8132 9234 8188
rect 9234 8132 9238 8188
rect 9174 8128 9238 8132
rect 9254 8188 9318 8192
rect 9254 8132 9258 8188
rect 9258 8132 9314 8188
rect 9314 8132 9318 8188
rect 9254 8128 9318 8132
rect 9334 8188 9398 8192
rect 9334 8132 9338 8188
rect 9338 8132 9394 8188
rect 9394 8132 9398 8188
rect 9334 8128 9398 8132
rect 14522 8188 14586 8192
rect 14522 8132 14526 8188
rect 14526 8132 14582 8188
rect 14582 8132 14586 8188
rect 14522 8128 14586 8132
rect 14602 8188 14666 8192
rect 14602 8132 14606 8188
rect 14606 8132 14662 8188
rect 14662 8132 14666 8188
rect 14602 8128 14666 8132
rect 14682 8188 14746 8192
rect 14682 8132 14686 8188
rect 14686 8132 14742 8188
rect 14742 8132 14746 8188
rect 14682 8128 14746 8132
rect 14762 8188 14826 8192
rect 14762 8132 14766 8188
rect 14766 8132 14822 8188
rect 14822 8132 14826 8188
rect 14762 8128 14826 8132
rect 19950 8188 20014 8192
rect 19950 8132 19954 8188
rect 19954 8132 20010 8188
rect 20010 8132 20014 8188
rect 19950 8128 20014 8132
rect 20030 8188 20094 8192
rect 20030 8132 20034 8188
rect 20034 8132 20090 8188
rect 20090 8132 20094 8188
rect 20030 8128 20094 8132
rect 20110 8188 20174 8192
rect 20110 8132 20114 8188
rect 20114 8132 20170 8188
rect 20170 8132 20174 8188
rect 20110 8128 20174 8132
rect 20190 8188 20254 8192
rect 20190 8132 20194 8188
rect 20194 8132 20250 8188
rect 20250 8132 20254 8188
rect 20190 8128 20254 8132
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 11808 7644 11872 7648
rect 11808 7588 11812 7644
rect 11812 7588 11868 7644
rect 11868 7588 11872 7644
rect 11808 7584 11872 7588
rect 11888 7644 11952 7648
rect 11888 7588 11892 7644
rect 11892 7588 11948 7644
rect 11948 7588 11952 7644
rect 11888 7584 11952 7588
rect 11968 7644 12032 7648
rect 11968 7588 11972 7644
rect 11972 7588 12028 7644
rect 12028 7588 12032 7644
rect 11968 7584 12032 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 17316 7644 17380 7648
rect 17316 7588 17320 7644
rect 17320 7588 17376 7644
rect 17376 7588 17380 7644
rect 17316 7584 17380 7588
rect 17396 7644 17460 7648
rect 17396 7588 17400 7644
rect 17400 7588 17456 7644
rect 17456 7588 17460 7644
rect 17396 7584 17460 7588
rect 17476 7644 17540 7648
rect 17476 7588 17480 7644
rect 17480 7588 17536 7644
rect 17536 7588 17540 7644
rect 17476 7584 17540 7588
rect 22664 7644 22728 7648
rect 22664 7588 22668 7644
rect 22668 7588 22724 7644
rect 22724 7588 22728 7644
rect 22664 7584 22728 7588
rect 22744 7644 22808 7648
rect 22744 7588 22748 7644
rect 22748 7588 22804 7644
rect 22804 7588 22808 7644
rect 22744 7584 22808 7588
rect 22824 7644 22888 7648
rect 22824 7588 22828 7644
rect 22828 7588 22884 7644
rect 22884 7588 22888 7644
rect 22824 7584 22888 7588
rect 22904 7644 22968 7648
rect 22904 7588 22908 7644
rect 22908 7588 22964 7644
rect 22964 7588 22968 7644
rect 22904 7584 22968 7588
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 9094 7100 9158 7104
rect 9094 7044 9098 7100
rect 9098 7044 9154 7100
rect 9154 7044 9158 7100
rect 9094 7040 9158 7044
rect 9174 7100 9238 7104
rect 9174 7044 9178 7100
rect 9178 7044 9234 7100
rect 9234 7044 9238 7100
rect 9174 7040 9238 7044
rect 9254 7100 9318 7104
rect 9254 7044 9258 7100
rect 9258 7044 9314 7100
rect 9314 7044 9318 7100
rect 9254 7040 9318 7044
rect 9334 7100 9398 7104
rect 9334 7044 9338 7100
rect 9338 7044 9394 7100
rect 9394 7044 9398 7100
rect 9334 7040 9398 7044
rect 14522 7100 14586 7104
rect 14522 7044 14526 7100
rect 14526 7044 14582 7100
rect 14582 7044 14586 7100
rect 14522 7040 14586 7044
rect 14602 7100 14666 7104
rect 14602 7044 14606 7100
rect 14606 7044 14662 7100
rect 14662 7044 14666 7100
rect 14602 7040 14666 7044
rect 14682 7100 14746 7104
rect 14682 7044 14686 7100
rect 14686 7044 14742 7100
rect 14742 7044 14746 7100
rect 14682 7040 14746 7044
rect 14762 7100 14826 7104
rect 14762 7044 14766 7100
rect 14766 7044 14822 7100
rect 14822 7044 14826 7100
rect 14762 7040 14826 7044
rect 19950 7100 20014 7104
rect 19950 7044 19954 7100
rect 19954 7044 20010 7100
rect 20010 7044 20014 7100
rect 19950 7040 20014 7044
rect 20030 7100 20094 7104
rect 20030 7044 20034 7100
rect 20034 7044 20090 7100
rect 20090 7044 20094 7100
rect 20030 7040 20094 7044
rect 20110 7100 20174 7104
rect 20110 7044 20114 7100
rect 20114 7044 20170 7100
rect 20170 7044 20174 7100
rect 20110 7040 20174 7044
rect 20190 7100 20254 7104
rect 20190 7044 20194 7100
rect 20194 7044 20250 7100
rect 20250 7044 20254 7100
rect 20190 7040 20254 7044
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 11808 6556 11872 6560
rect 11808 6500 11812 6556
rect 11812 6500 11868 6556
rect 11868 6500 11872 6556
rect 11808 6496 11872 6500
rect 11888 6556 11952 6560
rect 11888 6500 11892 6556
rect 11892 6500 11948 6556
rect 11948 6500 11952 6556
rect 11888 6496 11952 6500
rect 11968 6556 12032 6560
rect 11968 6500 11972 6556
rect 11972 6500 12028 6556
rect 12028 6500 12032 6556
rect 11968 6496 12032 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 17316 6556 17380 6560
rect 17316 6500 17320 6556
rect 17320 6500 17376 6556
rect 17376 6500 17380 6556
rect 17316 6496 17380 6500
rect 17396 6556 17460 6560
rect 17396 6500 17400 6556
rect 17400 6500 17456 6556
rect 17456 6500 17460 6556
rect 17396 6496 17460 6500
rect 17476 6556 17540 6560
rect 17476 6500 17480 6556
rect 17480 6500 17536 6556
rect 17536 6500 17540 6556
rect 17476 6496 17540 6500
rect 22664 6556 22728 6560
rect 22664 6500 22668 6556
rect 22668 6500 22724 6556
rect 22724 6500 22728 6556
rect 22664 6496 22728 6500
rect 22744 6556 22808 6560
rect 22744 6500 22748 6556
rect 22748 6500 22804 6556
rect 22804 6500 22808 6556
rect 22744 6496 22808 6500
rect 22824 6556 22888 6560
rect 22824 6500 22828 6556
rect 22828 6500 22884 6556
rect 22884 6500 22888 6556
rect 22824 6496 22888 6500
rect 22904 6556 22968 6560
rect 22904 6500 22908 6556
rect 22908 6500 22964 6556
rect 22964 6500 22968 6556
rect 22904 6496 22968 6500
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 9094 6012 9158 6016
rect 9094 5956 9098 6012
rect 9098 5956 9154 6012
rect 9154 5956 9158 6012
rect 9094 5952 9158 5956
rect 9174 6012 9238 6016
rect 9174 5956 9178 6012
rect 9178 5956 9234 6012
rect 9234 5956 9238 6012
rect 9174 5952 9238 5956
rect 9254 6012 9318 6016
rect 9254 5956 9258 6012
rect 9258 5956 9314 6012
rect 9314 5956 9318 6012
rect 9254 5952 9318 5956
rect 9334 6012 9398 6016
rect 9334 5956 9338 6012
rect 9338 5956 9394 6012
rect 9394 5956 9398 6012
rect 9334 5952 9398 5956
rect 14522 6012 14586 6016
rect 14522 5956 14526 6012
rect 14526 5956 14582 6012
rect 14582 5956 14586 6012
rect 14522 5952 14586 5956
rect 14602 6012 14666 6016
rect 14602 5956 14606 6012
rect 14606 5956 14662 6012
rect 14662 5956 14666 6012
rect 14602 5952 14666 5956
rect 14682 6012 14746 6016
rect 14682 5956 14686 6012
rect 14686 5956 14742 6012
rect 14742 5956 14746 6012
rect 14682 5952 14746 5956
rect 14762 6012 14826 6016
rect 14762 5956 14766 6012
rect 14766 5956 14822 6012
rect 14822 5956 14826 6012
rect 14762 5952 14826 5956
rect 19950 6012 20014 6016
rect 19950 5956 19954 6012
rect 19954 5956 20010 6012
rect 20010 5956 20014 6012
rect 19950 5952 20014 5956
rect 20030 6012 20094 6016
rect 20030 5956 20034 6012
rect 20034 5956 20090 6012
rect 20090 5956 20094 6012
rect 20030 5952 20094 5956
rect 20110 6012 20174 6016
rect 20110 5956 20114 6012
rect 20114 5956 20170 6012
rect 20170 5956 20174 6012
rect 20110 5952 20174 5956
rect 20190 6012 20254 6016
rect 20190 5956 20194 6012
rect 20194 5956 20250 6012
rect 20250 5956 20254 6012
rect 20190 5952 20254 5956
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 11808 5468 11872 5472
rect 11808 5412 11812 5468
rect 11812 5412 11868 5468
rect 11868 5412 11872 5468
rect 11808 5408 11872 5412
rect 11888 5468 11952 5472
rect 11888 5412 11892 5468
rect 11892 5412 11948 5468
rect 11948 5412 11952 5468
rect 11888 5408 11952 5412
rect 11968 5468 12032 5472
rect 11968 5412 11972 5468
rect 11972 5412 12028 5468
rect 12028 5412 12032 5468
rect 11968 5408 12032 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 17316 5468 17380 5472
rect 17316 5412 17320 5468
rect 17320 5412 17376 5468
rect 17376 5412 17380 5468
rect 17316 5408 17380 5412
rect 17396 5468 17460 5472
rect 17396 5412 17400 5468
rect 17400 5412 17456 5468
rect 17456 5412 17460 5468
rect 17396 5408 17460 5412
rect 17476 5468 17540 5472
rect 17476 5412 17480 5468
rect 17480 5412 17536 5468
rect 17536 5412 17540 5468
rect 17476 5408 17540 5412
rect 22664 5468 22728 5472
rect 22664 5412 22668 5468
rect 22668 5412 22724 5468
rect 22724 5412 22728 5468
rect 22664 5408 22728 5412
rect 22744 5468 22808 5472
rect 22744 5412 22748 5468
rect 22748 5412 22804 5468
rect 22804 5412 22808 5468
rect 22744 5408 22808 5412
rect 22824 5468 22888 5472
rect 22824 5412 22828 5468
rect 22828 5412 22884 5468
rect 22884 5412 22888 5468
rect 22824 5408 22888 5412
rect 22904 5468 22968 5472
rect 22904 5412 22908 5468
rect 22908 5412 22964 5468
rect 22964 5412 22968 5468
rect 22904 5408 22968 5412
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 9094 4924 9158 4928
rect 9094 4868 9098 4924
rect 9098 4868 9154 4924
rect 9154 4868 9158 4924
rect 9094 4864 9158 4868
rect 9174 4924 9238 4928
rect 9174 4868 9178 4924
rect 9178 4868 9234 4924
rect 9234 4868 9238 4924
rect 9174 4864 9238 4868
rect 9254 4924 9318 4928
rect 9254 4868 9258 4924
rect 9258 4868 9314 4924
rect 9314 4868 9318 4924
rect 9254 4864 9318 4868
rect 9334 4924 9398 4928
rect 9334 4868 9338 4924
rect 9338 4868 9394 4924
rect 9394 4868 9398 4924
rect 9334 4864 9398 4868
rect 14522 4924 14586 4928
rect 14522 4868 14526 4924
rect 14526 4868 14582 4924
rect 14582 4868 14586 4924
rect 14522 4864 14586 4868
rect 14602 4924 14666 4928
rect 14602 4868 14606 4924
rect 14606 4868 14662 4924
rect 14662 4868 14666 4924
rect 14602 4864 14666 4868
rect 14682 4924 14746 4928
rect 14682 4868 14686 4924
rect 14686 4868 14742 4924
rect 14742 4868 14746 4924
rect 14682 4864 14746 4868
rect 14762 4924 14826 4928
rect 14762 4868 14766 4924
rect 14766 4868 14822 4924
rect 14822 4868 14826 4924
rect 14762 4864 14826 4868
rect 19950 4924 20014 4928
rect 19950 4868 19954 4924
rect 19954 4868 20010 4924
rect 20010 4868 20014 4924
rect 19950 4864 20014 4868
rect 20030 4924 20094 4928
rect 20030 4868 20034 4924
rect 20034 4868 20090 4924
rect 20090 4868 20094 4924
rect 20030 4864 20094 4868
rect 20110 4924 20174 4928
rect 20110 4868 20114 4924
rect 20114 4868 20170 4924
rect 20170 4868 20174 4924
rect 20110 4864 20174 4868
rect 20190 4924 20254 4928
rect 20190 4868 20194 4924
rect 20194 4868 20250 4924
rect 20250 4868 20254 4924
rect 20190 4864 20254 4868
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 11808 4380 11872 4384
rect 11808 4324 11812 4380
rect 11812 4324 11868 4380
rect 11868 4324 11872 4380
rect 11808 4320 11872 4324
rect 11888 4380 11952 4384
rect 11888 4324 11892 4380
rect 11892 4324 11948 4380
rect 11948 4324 11952 4380
rect 11888 4320 11952 4324
rect 11968 4380 12032 4384
rect 11968 4324 11972 4380
rect 11972 4324 12028 4380
rect 12028 4324 12032 4380
rect 11968 4320 12032 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 17316 4380 17380 4384
rect 17316 4324 17320 4380
rect 17320 4324 17376 4380
rect 17376 4324 17380 4380
rect 17316 4320 17380 4324
rect 17396 4380 17460 4384
rect 17396 4324 17400 4380
rect 17400 4324 17456 4380
rect 17456 4324 17460 4380
rect 17396 4320 17460 4324
rect 17476 4380 17540 4384
rect 17476 4324 17480 4380
rect 17480 4324 17536 4380
rect 17536 4324 17540 4380
rect 17476 4320 17540 4324
rect 22664 4380 22728 4384
rect 22664 4324 22668 4380
rect 22668 4324 22724 4380
rect 22724 4324 22728 4380
rect 22664 4320 22728 4324
rect 22744 4380 22808 4384
rect 22744 4324 22748 4380
rect 22748 4324 22804 4380
rect 22804 4324 22808 4380
rect 22744 4320 22808 4324
rect 22824 4380 22888 4384
rect 22824 4324 22828 4380
rect 22828 4324 22884 4380
rect 22884 4324 22888 4380
rect 22824 4320 22888 4324
rect 22904 4380 22968 4384
rect 22904 4324 22908 4380
rect 22908 4324 22964 4380
rect 22964 4324 22968 4380
rect 22904 4320 22968 4324
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 9094 3836 9158 3840
rect 9094 3780 9098 3836
rect 9098 3780 9154 3836
rect 9154 3780 9158 3836
rect 9094 3776 9158 3780
rect 9174 3836 9238 3840
rect 9174 3780 9178 3836
rect 9178 3780 9234 3836
rect 9234 3780 9238 3836
rect 9174 3776 9238 3780
rect 9254 3836 9318 3840
rect 9254 3780 9258 3836
rect 9258 3780 9314 3836
rect 9314 3780 9318 3836
rect 9254 3776 9318 3780
rect 9334 3836 9398 3840
rect 9334 3780 9338 3836
rect 9338 3780 9394 3836
rect 9394 3780 9398 3836
rect 9334 3776 9398 3780
rect 14522 3836 14586 3840
rect 14522 3780 14526 3836
rect 14526 3780 14582 3836
rect 14582 3780 14586 3836
rect 14522 3776 14586 3780
rect 14602 3836 14666 3840
rect 14602 3780 14606 3836
rect 14606 3780 14662 3836
rect 14662 3780 14666 3836
rect 14602 3776 14666 3780
rect 14682 3836 14746 3840
rect 14682 3780 14686 3836
rect 14686 3780 14742 3836
rect 14742 3780 14746 3836
rect 14682 3776 14746 3780
rect 14762 3836 14826 3840
rect 14762 3780 14766 3836
rect 14766 3780 14822 3836
rect 14822 3780 14826 3836
rect 14762 3776 14826 3780
rect 19950 3836 20014 3840
rect 19950 3780 19954 3836
rect 19954 3780 20010 3836
rect 20010 3780 20014 3836
rect 19950 3776 20014 3780
rect 20030 3836 20094 3840
rect 20030 3780 20034 3836
rect 20034 3780 20090 3836
rect 20090 3780 20094 3836
rect 20030 3776 20094 3780
rect 20110 3836 20174 3840
rect 20110 3780 20114 3836
rect 20114 3780 20170 3836
rect 20170 3780 20174 3836
rect 20110 3776 20174 3780
rect 20190 3836 20254 3840
rect 20190 3780 20194 3836
rect 20194 3780 20250 3836
rect 20250 3780 20254 3836
rect 20190 3776 20254 3780
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 11808 3292 11872 3296
rect 11808 3236 11812 3292
rect 11812 3236 11868 3292
rect 11868 3236 11872 3292
rect 11808 3232 11872 3236
rect 11888 3292 11952 3296
rect 11888 3236 11892 3292
rect 11892 3236 11948 3292
rect 11948 3236 11952 3292
rect 11888 3232 11952 3236
rect 11968 3292 12032 3296
rect 11968 3236 11972 3292
rect 11972 3236 12028 3292
rect 12028 3236 12032 3292
rect 11968 3232 12032 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 17316 3292 17380 3296
rect 17316 3236 17320 3292
rect 17320 3236 17376 3292
rect 17376 3236 17380 3292
rect 17316 3232 17380 3236
rect 17396 3292 17460 3296
rect 17396 3236 17400 3292
rect 17400 3236 17456 3292
rect 17456 3236 17460 3292
rect 17396 3232 17460 3236
rect 17476 3292 17540 3296
rect 17476 3236 17480 3292
rect 17480 3236 17536 3292
rect 17536 3236 17540 3292
rect 17476 3232 17540 3236
rect 22664 3292 22728 3296
rect 22664 3236 22668 3292
rect 22668 3236 22724 3292
rect 22724 3236 22728 3292
rect 22664 3232 22728 3236
rect 22744 3292 22808 3296
rect 22744 3236 22748 3292
rect 22748 3236 22804 3292
rect 22804 3236 22808 3292
rect 22744 3232 22808 3236
rect 22824 3292 22888 3296
rect 22824 3236 22828 3292
rect 22828 3236 22884 3292
rect 22884 3236 22888 3292
rect 22824 3232 22888 3236
rect 22904 3292 22968 3296
rect 22904 3236 22908 3292
rect 22908 3236 22964 3292
rect 22964 3236 22968 3292
rect 22904 3232 22968 3236
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 9094 2748 9158 2752
rect 9094 2692 9098 2748
rect 9098 2692 9154 2748
rect 9154 2692 9158 2748
rect 9094 2688 9158 2692
rect 9174 2748 9238 2752
rect 9174 2692 9178 2748
rect 9178 2692 9234 2748
rect 9234 2692 9238 2748
rect 9174 2688 9238 2692
rect 9254 2748 9318 2752
rect 9254 2692 9258 2748
rect 9258 2692 9314 2748
rect 9314 2692 9318 2748
rect 9254 2688 9318 2692
rect 9334 2748 9398 2752
rect 9334 2692 9338 2748
rect 9338 2692 9394 2748
rect 9394 2692 9398 2748
rect 9334 2688 9398 2692
rect 14522 2748 14586 2752
rect 14522 2692 14526 2748
rect 14526 2692 14582 2748
rect 14582 2692 14586 2748
rect 14522 2688 14586 2692
rect 14602 2748 14666 2752
rect 14602 2692 14606 2748
rect 14606 2692 14662 2748
rect 14662 2692 14666 2748
rect 14602 2688 14666 2692
rect 14682 2748 14746 2752
rect 14682 2692 14686 2748
rect 14686 2692 14742 2748
rect 14742 2692 14746 2748
rect 14682 2688 14746 2692
rect 14762 2748 14826 2752
rect 14762 2692 14766 2748
rect 14766 2692 14822 2748
rect 14822 2692 14826 2748
rect 14762 2688 14826 2692
rect 19950 2748 20014 2752
rect 19950 2692 19954 2748
rect 19954 2692 20010 2748
rect 20010 2692 20014 2748
rect 19950 2688 20014 2692
rect 20030 2748 20094 2752
rect 20030 2692 20034 2748
rect 20034 2692 20090 2748
rect 20090 2692 20094 2748
rect 20030 2688 20094 2692
rect 20110 2748 20174 2752
rect 20110 2692 20114 2748
rect 20114 2692 20170 2748
rect 20170 2692 20174 2748
rect 20110 2688 20174 2692
rect 20190 2748 20254 2752
rect 20190 2692 20194 2748
rect 20194 2692 20250 2748
rect 20250 2692 20254 2748
rect 20190 2688 20254 2692
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 11808 2204 11872 2208
rect 11808 2148 11812 2204
rect 11812 2148 11868 2204
rect 11868 2148 11872 2204
rect 11808 2144 11872 2148
rect 11888 2204 11952 2208
rect 11888 2148 11892 2204
rect 11892 2148 11948 2204
rect 11948 2148 11952 2204
rect 11888 2144 11952 2148
rect 11968 2204 12032 2208
rect 11968 2148 11972 2204
rect 11972 2148 12028 2204
rect 12028 2148 12032 2204
rect 11968 2144 12032 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 17316 2204 17380 2208
rect 17316 2148 17320 2204
rect 17320 2148 17376 2204
rect 17376 2148 17380 2204
rect 17316 2144 17380 2148
rect 17396 2204 17460 2208
rect 17396 2148 17400 2204
rect 17400 2148 17456 2204
rect 17456 2148 17460 2204
rect 17396 2144 17460 2148
rect 17476 2204 17540 2208
rect 17476 2148 17480 2204
rect 17480 2148 17536 2204
rect 17536 2148 17540 2204
rect 17476 2144 17540 2148
rect 22664 2204 22728 2208
rect 22664 2148 22668 2204
rect 22668 2148 22724 2204
rect 22724 2148 22728 2204
rect 22664 2144 22728 2148
rect 22744 2204 22808 2208
rect 22744 2148 22748 2204
rect 22748 2148 22804 2204
rect 22804 2148 22808 2204
rect 22744 2144 22808 2148
rect 22824 2204 22888 2208
rect 22824 2148 22828 2204
rect 22828 2148 22884 2204
rect 22884 2148 22888 2204
rect 22824 2144 22888 2148
rect 22904 2204 22968 2208
rect 22904 2148 22908 2204
rect 22908 2148 22964 2204
rect 22964 2148 22968 2204
rect 22904 2144 22968 2148
<< metal4 >>
rect 3658 21248 3978 21808
rect 3658 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3978 21248
rect 3658 20160 3978 21184
rect 3658 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3978 20160
rect 3658 19072 3978 20096
rect 3658 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3978 19072
rect 3658 17984 3978 19008
rect 3658 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3978 17984
rect 3658 16896 3978 17920
rect 3658 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3978 16896
rect 3658 15808 3978 16832
rect 3658 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3978 15808
rect 3658 14720 3978 15744
rect 3658 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3978 14720
rect 3658 13632 3978 14656
rect 3658 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3978 13632
rect 3658 12544 3978 13568
rect 3658 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3978 12544
rect 3658 11456 3978 12480
rect 3658 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3978 11456
rect 3658 10368 3978 11392
rect 3658 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3978 10368
rect 3658 9280 3978 10304
rect 3658 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3978 9280
rect 3658 8192 3978 9216
rect 3658 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3978 8192
rect 3658 7104 3978 8128
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6016 3978 7040
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4928 3978 5952
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 3840 3978 4864
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 2752 3978 3776
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 6372 21792 6692 21808
rect 6372 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6692 21792
rect 6372 20704 6692 21728
rect 6372 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6692 20704
rect 6372 19616 6692 20640
rect 6372 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6692 19616
rect 6372 18528 6692 19552
rect 6372 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6692 18528
rect 6372 17440 6692 18464
rect 6372 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6692 17440
rect 6372 16352 6692 17376
rect 6372 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6692 16352
rect 6372 15264 6692 16288
rect 6372 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6692 15264
rect 6372 14176 6692 15200
rect 6372 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6692 14176
rect 6372 13088 6692 14112
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 10912 6692 11936
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7648 6692 8672
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 6560 6692 7584
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 5472 6692 6496
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 3296 6692 4320
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 9086 21248 9406 21808
rect 9086 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9406 21248
rect 9086 20160 9406 21184
rect 9086 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9406 20160
rect 9086 19072 9406 20096
rect 9086 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9406 19072
rect 9086 17984 9406 19008
rect 9086 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9406 17984
rect 9086 16896 9406 17920
rect 9086 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9406 16896
rect 9086 15808 9406 16832
rect 9086 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9406 15808
rect 9086 14720 9406 15744
rect 9086 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9406 14720
rect 9086 13632 9406 14656
rect 9086 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9406 13632
rect 9086 12544 9406 13568
rect 9086 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9406 12544
rect 9086 11456 9406 12480
rect 9086 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9406 11456
rect 9086 10368 9406 11392
rect 9086 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9406 10368
rect 9086 9280 9406 10304
rect 9086 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9406 9280
rect 9086 8192 9406 9216
rect 9086 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9406 8192
rect 9086 7104 9406 8128
rect 9086 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9406 7104
rect 9086 6016 9406 7040
rect 9086 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9406 6016
rect 9086 4928 9406 5952
rect 9086 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9406 4928
rect 9086 3840 9406 4864
rect 9086 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9406 3840
rect 9086 2752 9406 3776
rect 9086 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9406 2752
rect 9086 2128 9406 2688
rect 11800 21792 12120 21808
rect 11800 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12120 21792
rect 11800 20704 12120 21728
rect 11800 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12120 20704
rect 11800 19616 12120 20640
rect 11800 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12120 19616
rect 11800 18528 12120 19552
rect 11800 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12120 18528
rect 11800 17440 12120 18464
rect 11800 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12120 17440
rect 11800 16352 12120 17376
rect 11800 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12120 16352
rect 11800 15264 12120 16288
rect 11800 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12120 15264
rect 11800 14176 12120 15200
rect 11800 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12120 14176
rect 11800 13088 12120 14112
rect 11800 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12120 13088
rect 11800 12000 12120 13024
rect 11800 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12120 12000
rect 11800 10912 12120 11936
rect 11800 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12120 10912
rect 11800 9824 12120 10848
rect 11800 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12120 9824
rect 11800 8736 12120 9760
rect 11800 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12120 8736
rect 11800 7648 12120 8672
rect 11800 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12120 7648
rect 11800 6560 12120 7584
rect 11800 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12120 6560
rect 11800 5472 12120 6496
rect 11800 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12120 5472
rect 11800 4384 12120 5408
rect 11800 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12120 4384
rect 11800 3296 12120 4320
rect 11800 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12120 3296
rect 11800 2208 12120 3232
rect 11800 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12120 2208
rect 11800 2128 12120 2144
rect 14514 21248 14834 21808
rect 14514 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14834 21248
rect 14514 20160 14834 21184
rect 14514 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14834 20160
rect 14514 19072 14834 20096
rect 14514 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14834 19072
rect 14514 17984 14834 19008
rect 14514 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14834 17984
rect 14514 16896 14834 17920
rect 14514 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14834 16896
rect 14514 15808 14834 16832
rect 14514 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14834 15808
rect 14514 14720 14834 15744
rect 14514 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14834 14720
rect 14514 13632 14834 14656
rect 14514 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14834 13632
rect 14514 12544 14834 13568
rect 14514 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14834 12544
rect 14514 11456 14834 12480
rect 14514 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14834 11456
rect 14514 10368 14834 11392
rect 14514 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14834 10368
rect 14514 9280 14834 10304
rect 14514 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14834 9280
rect 14514 8192 14834 9216
rect 14514 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14834 8192
rect 14514 7104 14834 8128
rect 14514 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14834 7104
rect 14514 6016 14834 7040
rect 14514 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14834 6016
rect 14514 4928 14834 5952
rect 14514 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14834 4928
rect 14514 3840 14834 4864
rect 14514 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14834 3840
rect 14514 2752 14834 3776
rect 14514 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14834 2752
rect 14514 2128 14834 2688
rect 17228 21792 17548 21808
rect 17228 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17548 21792
rect 17228 20704 17548 21728
rect 17228 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17548 20704
rect 17228 19616 17548 20640
rect 17228 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17548 19616
rect 17228 18528 17548 19552
rect 17228 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17548 18528
rect 17228 17440 17548 18464
rect 17228 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17548 17440
rect 17228 16352 17548 17376
rect 17228 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17548 16352
rect 17228 15264 17548 16288
rect 17228 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17548 15264
rect 17228 14176 17548 15200
rect 17228 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17548 14176
rect 17228 13088 17548 14112
rect 17228 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17548 13088
rect 17228 12000 17548 13024
rect 17228 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17548 12000
rect 17228 10912 17548 11936
rect 17228 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17548 10912
rect 17228 9824 17548 10848
rect 17228 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17548 9824
rect 17228 8736 17548 9760
rect 17228 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17548 8736
rect 17228 7648 17548 8672
rect 17228 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17548 7648
rect 17228 6560 17548 7584
rect 17228 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17548 6560
rect 17228 5472 17548 6496
rect 17228 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17548 5472
rect 17228 4384 17548 5408
rect 17228 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17548 4384
rect 17228 3296 17548 4320
rect 17228 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17548 3296
rect 17228 2208 17548 3232
rect 17228 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17548 2208
rect 17228 2128 17548 2144
rect 19942 21248 20262 21808
rect 19942 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20262 21248
rect 19942 20160 20262 21184
rect 19942 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20262 20160
rect 19942 19072 20262 20096
rect 19942 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20262 19072
rect 19942 17984 20262 19008
rect 19942 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20262 17984
rect 19942 16896 20262 17920
rect 19942 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20262 16896
rect 19942 15808 20262 16832
rect 19942 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20262 15808
rect 19942 14720 20262 15744
rect 19942 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20262 14720
rect 19942 13632 20262 14656
rect 19942 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20262 13632
rect 19942 12544 20262 13568
rect 19942 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20262 12544
rect 19942 11456 20262 12480
rect 19942 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20262 11456
rect 19942 10368 20262 11392
rect 19942 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20262 10368
rect 19942 9280 20262 10304
rect 19942 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20262 9280
rect 19942 8192 20262 9216
rect 19942 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20262 8192
rect 19942 7104 20262 8128
rect 19942 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20262 7104
rect 19942 6016 20262 7040
rect 19942 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20262 6016
rect 19942 4928 20262 5952
rect 19942 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20262 4928
rect 19942 3840 20262 4864
rect 19942 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20262 3840
rect 19942 2752 20262 3776
rect 19942 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20262 2752
rect 19942 2128 20262 2688
rect 22656 21792 22976 21808
rect 22656 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22976 21792
rect 22656 20704 22976 21728
rect 22656 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22976 20704
rect 22656 19616 22976 20640
rect 22656 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22976 19616
rect 22656 18528 22976 19552
rect 22656 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22976 18528
rect 22656 17440 22976 18464
rect 22656 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22976 17440
rect 22656 16352 22976 17376
rect 22656 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22976 16352
rect 22656 15264 22976 16288
rect 22656 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22976 15264
rect 22656 14176 22976 15200
rect 22656 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22976 14176
rect 22656 13088 22976 14112
rect 22656 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22976 13088
rect 22656 12000 22976 13024
rect 22656 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22976 12000
rect 22656 10912 22976 11936
rect 22656 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22976 10912
rect 22656 9824 22976 10848
rect 22656 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22976 9824
rect 22656 8736 22976 9760
rect 22656 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22976 8736
rect 22656 7648 22976 8672
rect 22656 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22976 7648
rect 22656 6560 22976 7584
rect 22656 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22976 6560
rect 22656 5472 22976 6496
rect 22656 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22976 5472
rect 22656 4384 22976 5408
rect 22656 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22976 4384
rect 22656 3296 22976 4320
rect 22656 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22976 3296
rect 22656 2208 22976 3232
rect 22656 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22976 2208
rect 22656 2128 22976 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A0 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20240 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A1
timestamp 1666464484
transform -1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A2
timestamp 1666464484
transform -1 0 18308 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A3
timestamp 1666464484
transform -1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_reg_clk_A
timestamp 1666464484
transform -1 0 22356 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 7360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 10856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 15088 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output6_A
timestamp 1666464484
transform 1 0 5428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output7_A
timestamp 1666464484
transform 1 0 8372 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_A
timestamp 1666464484
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp 1666464484
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1666464484
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68
timestamp 1666464484
transform 1 0 7360 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1666464484
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1666464484
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1666464484
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152
timestamp 1666464484
transform 1 0 15088 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1666464484
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1666464484
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_230
timestamp 1666464484
transform 1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1666464484
transform 1 0 14628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1666464484
transform 1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1666464484
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1666464484
transform 1 0 17112 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_203
timestamp 1666464484
transform 1 0 19780 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1666464484
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_230
timestamp 1666464484
transform 1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1666464484
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_231
timestamp 1666464484
transform 1 0 22356 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_197
timestamp 1666464484
transform 1 0 19228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1666464484
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_230
timestamp 1666464484
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_185
timestamp 1666464484
transform 1 0 18124 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666464484
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1666464484
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_206
timestamp 1666464484
transform 1 0 20056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1666464484
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_228
timestamp 1666464484
transform 1 0 22080 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_231
timestamp 1666464484
transform 1 0 22356 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_206
timestamp 1666464484
transform 1 0 20056 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_210
timestamp 1666464484
transform 1 0 20424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 1666464484
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1666464484
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_205
timestamp 1666464484
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_222
timestamp 1666464484
transform 1 0 21528 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_230
timestamp 1666464484
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1666464484
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1666464484
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_194
timestamp 1666464484
transform 1 0 18952 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_206
timestamp 1666464484
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1666464484
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_183
timestamp 1666464484
transform 1 0 17940 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_204
timestamp 1666464484
transform 1 0 19872 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_216
timestamp 1666464484
transform 1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_228
timestamp 1666464484
transform 1 0 22080 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_232
timestamp 1666464484
transform 1 0 22448 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_189
timestamp 1666464484
transform 1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_197
timestamp 1666464484
transform 1 0 19228 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_212
timestamp 1666464484
transform 1 0 20608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1666464484
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_231
timestamp 1666464484
transform 1 0 22356 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1666464484
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1666464484
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1666464484
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_207
timestamp 1666464484
transform 1 0 20148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_215
timestamp 1666464484
transform 1 0 20884 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1666464484
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1666464484
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1666464484
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_211
timestamp 1666464484
transform 1 0 20516 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_229
timestamp 1666464484
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_183
timestamp 1666464484
transform 1 0 17940 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1666464484
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1666464484
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_208
timestamp 1666464484
transform 1 0 20240 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1666464484
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_173
timestamp 1666464484
transform 1 0 17020 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_184
timestamp 1666464484
transform 1 0 18032 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1666464484
transform 1 0 18032 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_194
timestamp 1666464484
transform 1 0 18952 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_206
timestamp 1666464484
transform 1 0 20056 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1666464484
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1666464484
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_175
timestamp 1666464484
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_211
timestamp 1666464484
transform 1 0 20516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_223
timestamp 1666464484
transform 1 0 21620 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1666464484
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_174
timestamp 1666464484
transform 1 0 17112 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_182
timestamp 1666464484
transform 1 0 17848 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_206
timestamp 1666464484
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1666464484
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_181
timestamp 1666464484
transform 1 0 17756 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1666464484
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_183
timestamp 1666464484
transform 1 0 17940 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_195
timestamp 1666464484
transform 1 0 19044 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_207
timestamp 1666464484
transform 1 0 20148 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1666464484
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_11
timestamp 1666464484
transform 1 0 2116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_17
timestamp 1666464484
transform 1 0 2668 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_25
timestamp 1666464484
transform 1 0 3404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_29
timestamp 1666464484
transform 1 0 3772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_37
timestamp 1666464484
transform 1 0 4508 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_43
timestamp 1666464484
transform 1 0 5060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_49
timestamp 1666464484
transform 1 0 5612 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1666464484
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_85
timestamp 1666464484
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_97
timestamp 1666464484
transform 1 0 10028 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1666464484
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_117
timestamp 1666464484
transform 1 0 11868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_129
timestamp 1666464484
transform 1 0 12972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_141
timestamp 1666464484
transform 1 0 14076 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_147
timestamp 1666464484
transform 1 0 14628 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1666464484
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_175
timestamp 1666464484
transform 1 0 17204 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_187
timestamp 1666464484
transform 1 0 18308 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_195
timestamp 1666464484
transform 1 0 19044 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1666464484
transform 1 0 19228 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_203
timestamp 1666464484
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_215
timestamp 1666464484
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_231
timestamp 1666464484
transform 1 0 22356 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 22816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 22816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 22816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _34_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20976 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _35_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21252 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _36_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _37_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20976 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _38_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20976 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _39_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _40_
timestamp 1666464484
transform -1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1666464484
transform -1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _43_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12972 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_2  _44_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _45_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _46_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18952 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _47_
timestamp 1666464484
transform 1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _48_
timestamp 1666464484
transform -1 0 18952 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _49_
timestamp 1666464484
transform -1 0 16376 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _50_
timestamp 1666464484
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _51_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18952 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _52_
timestamp 1666464484
transform 1 0 17112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _53_
timestamp 1666464484
transform -1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _54_
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _55_
timestamp 1666464484
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _56__1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19320 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _57__2
timestamp 1666464484
transform 1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _58__3
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _59__4
timestamp 1666464484
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _60_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20056 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _61_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _62_
timestamp 1666464484
transform 1 0 17020 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _63_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19228 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _64_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14076 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _65_
timestamp 1666464484
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _66_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18952 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _67_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _68_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _69_
timestamp 1666464484
transform -1 0 18952 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _70_
timestamp 1666464484
transform -1 0 21712 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _70__13 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _71_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _72_
timestamp 1666464484
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _73_
timestamp 1666464484
transform 1 0 16652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _74_
timestamp 1666464484
transform 1 0 18584 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _75_
timestamp 1666464484
transform 1 0 16928 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _76_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _77_
timestamp 1666464484
transform 1 0 19412 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _78_
timestamp 1666464484
transform 1 0 19412 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _79_
timestamp 1666464484
transform 1 0 20056 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__ebufn_8  _81_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17848 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_reg_clk dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22356 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_reg_clk
timestamp 1666464484
transform 1 0 19688 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_reg_clk
timestamp 1666464484
transform -1 0 20056 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform -1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output5 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform -1 0 5060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform -1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform -1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform -1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform -1 0 19780 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform 1 0 21988 0 -1 21760
box -38 -48 406 592
<< labels >>
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 reg_addr[0]
port 0 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 reg_addr[1]
port 1 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 reg_addr[2]
port 2 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 reg_bus
port 3 nsew signal bidirectional
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 reg_clk
port 4 nsew signal input
flabel metal2 s 1674 23200 1730 24000 0 FreeSans 224 90 0 0 reg_data[0]
port 5 nsew signal tristate
flabel metal2 s 4618 23200 4674 24000 0 FreeSans 224 90 0 0 reg_data[1]
port 6 nsew signal tristate
flabel metal2 s 7562 23200 7618 24000 0 FreeSans 224 90 0 0 reg_data[2]
port 7 nsew signal tristate
flabel metal2 s 10506 23200 10562 24000 0 FreeSans 224 90 0 0 reg_data[3]
port 8 nsew signal tristate
flabel metal2 s 13450 23200 13506 24000 0 FreeSans 224 90 0 0 reg_data[4]
port 9 nsew signal tristate
flabel metal2 s 16394 23200 16450 24000 0 FreeSans 224 90 0 0 reg_data[5]
port 10 nsew signal tristate
flabel metal2 s 19338 23200 19394 24000 0 FreeSans 224 90 0 0 reg_data[6]
port 11 nsew signal tristate
flabel metal2 s 22282 23200 22338 24000 0 FreeSans 224 90 0 0 reg_data[7]
port 12 nsew signal tristate
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 reg_dir
port 13 nsew signal input
flabel metal4 s 3658 2128 3978 21808 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 9086 2128 9406 21808 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 14514 2128 14834 21808 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 19942 2128 20262 21808 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 6372 2128 6692 21808 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 11800 2128 12120 21808 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 17228 2128 17548 21808 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 22656 2128 22976 21808 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
rlabel metal1 11960 21216 11960 21216 0 vccd1
rlabel via1 12040 21760 12040 21760 0 vssd1
rlabel metal2 17894 10812 17894 10812 0 _00_
rlabel metal1 15870 12274 15870 12274 0 _01_
rlabel metal2 16238 13124 16238 13124 0 _02_
rlabel metal1 18722 9690 18722 9690 0 _03_
rlabel metal2 16974 11492 16974 11492 0 _04_
rlabel metal2 16882 13396 16882 13396 0 _05_
rlabel metal1 19090 13158 19090 13158 0 _06_
rlabel metal2 19458 9860 19458 9860 0 _07_
rlabel metal1 18952 3706 18952 3706 0 _12_
rlabel metal1 20419 6358 20419 6358 0 _13_
rlabel metal1 19841 2346 19841 2346 0 _14_
rlabel metal1 19274 4794 19274 4794 0 _16_
rlabel metal2 21298 10268 21298 10268 0 _17_
rlabel metal1 17572 11118 17572 11118 0 _18_
rlabel metal1 21620 8330 21620 8330 0 _19_
rlabel metal1 19550 9520 19550 9520 0 _20_
rlabel metal1 16330 3026 16330 3026 0 _21_
rlabel metal2 18446 5236 18446 5236 0 _22_
rlabel metal2 18722 8670 18722 8670 0 _23_
rlabel metal1 17664 11526 17664 11526 0 _24_
rlabel metal1 18262 12648 18262 12648 0 _25_
rlabel metal1 17526 12818 17526 12818 0 _26_
rlabel metal1 18814 7922 18814 7922 0 _27_
rlabel metal2 18538 6120 18538 6120 0 _28_
rlabel metal2 18906 9078 18906 9078 0 _29_
rlabel metal2 18630 6460 18630 6460 0 _30_
rlabel metal1 19458 4624 19458 4624 0 _31_
rlabel metal1 18722 4556 18722 4556 0 _32_
rlabel metal1 18078 2924 18078 2924 0 _33_
rlabel metal1 20286 2414 20286 2414 0 clknet_0_reg_clk
rlabel metal1 21758 2414 21758 2414 0 clknet_1_0__leaf_reg_clk
rlabel metal2 19366 4556 19366 4556 0 clknet_1_1__leaf_reg_clk
rlabel metal2 18262 5100 18262 5100 0 data_t
rlabel metal1 10074 2278 10074 2278 0 net1
rlabel metal1 17526 21522 17526 21522 0 net10
rlabel metal1 20102 21522 20102 21522 0 net11
rlabel metal1 20930 21454 20930 21454 0 net12
rlabel metal2 22034 4318 22034 4318 0 net13
rlabel metal1 19734 4046 19734 4046 0 net14
rlabel metal1 20562 5338 20562 5338 0 net15
rlabel metal1 20516 2482 20516 2482 0 net16
rlabel metal2 22126 3876 22126 3876 0 net17
rlabel metal2 12374 2788 12374 2788 0 net2
rlabel metal1 14214 2618 14214 2618 0 net3
rlabel metal1 7682 2550 7682 2550 0 net4
rlabel metal1 2300 21522 2300 21522 0 net5
rlabel metal1 5888 21318 5888 21318 0 net6
rlabel metal1 8188 21522 8188 21522 0 net7
rlabel metal1 11316 21522 11316 21522 0 net8
rlabel metal2 19090 17136 19090 17136 0 net9
rlabel metal1 6302 2414 6302 2414 0 reg_addr[0]
rlabel metal1 10028 2414 10028 2414 0 reg_addr[1]
rlabel metal1 14214 2414 14214 2414 0 reg_addr[2]
rlabel metal1 17112 13906 17112 13906 0 reg_bus
rlabel metal2 22218 3944 22218 3944 0 reg_clk
rlabel metal2 1886 22491 1886 22491 0 reg_data[0]
rlabel metal2 4830 22491 4830 22491 0 reg_data[1]
rlabel metal2 7774 22491 7774 22491 0 reg_data[2]
rlabel metal2 10718 22491 10718 22491 0 reg_data[3]
rlabel metal1 14122 21658 14122 21658 0 reg_data[4]
rlabel metal1 16790 21658 16790 21658 0 reg_data[5]
rlabel metal2 19550 22491 19550 22491 0 reg_data[6]
rlabel metal2 22218 22491 22218 22491 0 reg_data[7]
rlabel metal1 2116 2414 2116 2414 0 reg_dir
rlabel metal1 19366 12648 19366 12648 0 t\[0\]
rlabel metal2 21206 7990 21206 7990 0 t\[1\]
rlabel metal1 18216 2618 18216 2618 0 t\[2\]
rlabel metal2 20562 8602 20562 8602 0 t\[3\]
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
