magic
tech sky130A
magscale 1 2
timestamp 1673257823
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 212 178848 117552
<< metal2 >>
rect 1582 119200 1638 120000
rect 3146 119200 3202 120000
rect 4710 119200 4766 120000
rect 6274 119200 6330 120000
rect 7838 119200 7894 120000
rect 9402 119200 9458 120000
rect 10966 119200 11022 120000
rect 12530 119200 12586 120000
rect 14094 119200 14150 120000
rect 15658 119200 15714 120000
rect 17222 119200 17278 120000
rect 18786 119200 18842 120000
rect 20350 119200 20406 120000
rect 21914 119200 21970 120000
rect 23478 119200 23534 120000
rect 25042 119200 25098 120000
rect 26606 119200 26662 120000
rect 28170 119200 28226 120000
rect 29734 119200 29790 120000
rect 31298 119200 31354 120000
rect 32862 119200 32918 120000
rect 34426 119200 34482 120000
rect 35990 119200 36046 120000
rect 37554 119200 37610 120000
rect 39118 119200 39174 120000
rect 40682 119200 40738 120000
rect 42246 119200 42302 120000
rect 43810 119200 43866 120000
rect 45374 119200 45430 120000
rect 46938 119200 46994 120000
rect 48502 119200 48558 120000
rect 50066 119200 50122 120000
rect 51630 119200 51686 120000
rect 53194 119200 53250 120000
rect 54758 119200 54814 120000
rect 56322 119200 56378 120000
rect 57886 119200 57942 120000
rect 59450 119200 59506 120000
rect 61014 119200 61070 120000
rect 62578 119200 62634 120000
rect 64142 119200 64198 120000
rect 65706 119200 65762 120000
rect 67270 119200 67326 120000
rect 68834 119200 68890 120000
rect 70398 119200 70454 120000
rect 71962 119200 72018 120000
rect 73526 119200 73582 120000
rect 75090 119200 75146 120000
rect 76654 119200 76710 120000
rect 78218 119200 78274 120000
rect 79782 119200 79838 120000
rect 81346 119200 81402 120000
rect 82910 119200 82966 120000
rect 84474 119200 84530 120000
rect 86038 119200 86094 120000
rect 87602 119200 87658 120000
rect 89166 119200 89222 120000
rect 90730 119200 90786 120000
rect 92294 119200 92350 120000
rect 93858 119200 93914 120000
rect 95422 119200 95478 120000
rect 96986 119200 97042 120000
rect 98550 119200 98606 120000
rect 100114 119200 100170 120000
rect 101678 119200 101734 120000
rect 103242 119200 103298 120000
rect 104806 119200 104862 120000
rect 106370 119200 106426 120000
rect 107934 119200 107990 120000
rect 109498 119200 109554 120000
rect 111062 119200 111118 120000
rect 112626 119200 112682 120000
rect 114190 119200 114246 120000
rect 115754 119200 115810 120000
rect 117318 119200 117374 120000
rect 118882 119200 118938 120000
rect 120446 119200 120502 120000
rect 122010 119200 122066 120000
rect 123574 119200 123630 120000
rect 125138 119200 125194 120000
rect 126702 119200 126758 120000
rect 128266 119200 128322 120000
rect 129830 119200 129886 120000
rect 131394 119200 131450 120000
rect 132958 119200 133014 120000
rect 134522 119200 134578 120000
rect 136086 119200 136142 120000
rect 137650 119200 137706 120000
rect 139214 119200 139270 120000
rect 140778 119200 140834 120000
rect 142342 119200 142398 120000
rect 143906 119200 143962 120000
rect 145470 119200 145526 120000
rect 147034 119200 147090 120000
rect 148598 119200 148654 120000
rect 150162 119200 150218 120000
rect 151726 119200 151782 120000
rect 153290 119200 153346 120000
rect 154854 119200 154910 120000
rect 156418 119200 156474 120000
rect 157982 119200 158038 120000
rect 159546 119200 159602 120000
rect 161110 119200 161166 120000
rect 162674 119200 162730 120000
rect 164238 119200 164294 120000
rect 165802 119200 165858 120000
rect 167366 119200 167422 120000
rect 168930 119200 168986 120000
rect 170494 119200 170550 120000
rect 172058 119200 172114 120000
rect 173622 119200 173678 120000
rect 175186 119200 175242 120000
rect 176750 119200 176806 120000
rect 178314 119200 178370 120000
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8206 0 8262 800
rect 8758 0 8814 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10414 0 10470 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17590 0 17646 800
rect 18142 0 18198 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23662 0 23718 800
rect 24214 0 24270 800
rect 24766 0 24822 800
rect 25318 0 25374 800
rect 25870 0 25926 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27526 0 27582 800
rect 28078 0 28134 800
rect 28630 0 28686 800
rect 29182 0 29238 800
rect 29734 0 29790 800
rect 30286 0 30342 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40222 0 40278 800
rect 40774 0 40830 800
rect 41326 0 41382 800
rect 41878 0 41934 800
rect 42430 0 42486 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44638 0 44694 800
rect 45190 0 45246 800
rect 45742 0 45798 800
rect 46294 0 46350 800
rect 46846 0 46902 800
rect 47398 0 47454 800
rect 47950 0 48006 800
rect 48502 0 48558 800
rect 49054 0 49110 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51262 0 51318 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52918 0 52974 800
rect 53470 0 53526 800
rect 54022 0 54078 800
rect 54574 0 54630 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56230 0 56286 800
rect 56782 0 56838 800
rect 57334 0 57390 800
rect 57886 0 57942 800
rect 58438 0 58494 800
rect 58990 0 59046 800
rect 59542 0 59598 800
rect 60094 0 60150 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64510 0 64566 800
rect 65062 0 65118 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66718 0 66774 800
rect 67270 0 67326 800
rect 67822 0 67878 800
rect 68374 0 68430 800
rect 68926 0 68982 800
rect 69478 0 69534 800
rect 70030 0 70086 800
rect 70582 0 70638 800
rect 71134 0 71190 800
rect 71686 0 71742 800
rect 72238 0 72294 800
rect 72790 0 72846 800
rect 73342 0 73398 800
rect 73894 0 73950 800
rect 74446 0 74502 800
rect 74998 0 75054 800
rect 75550 0 75606 800
rect 76102 0 76158 800
rect 76654 0 76710 800
rect 77206 0 77262 800
rect 77758 0 77814 800
rect 78310 0 78366 800
rect 78862 0 78918 800
rect 79414 0 79470 800
rect 79966 0 80022 800
rect 80518 0 80574 800
rect 81070 0 81126 800
rect 81622 0 81678 800
rect 82174 0 82230 800
rect 82726 0 82782 800
rect 83278 0 83334 800
rect 83830 0 83886 800
rect 84382 0 84438 800
rect 84934 0 84990 800
rect 85486 0 85542 800
rect 86038 0 86094 800
rect 86590 0 86646 800
rect 87142 0 87198 800
rect 87694 0 87750 800
rect 88246 0 88302 800
rect 88798 0 88854 800
rect 89350 0 89406 800
rect 89902 0 89958 800
rect 90454 0 90510 800
rect 91006 0 91062 800
rect 91558 0 91614 800
rect 92110 0 92166 800
rect 92662 0 92718 800
rect 93214 0 93270 800
rect 93766 0 93822 800
rect 94318 0 94374 800
rect 94870 0 94926 800
rect 95422 0 95478 800
rect 95974 0 96030 800
rect 96526 0 96582 800
rect 97078 0 97134 800
rect 97630 0 97686 800
rect 98182 0 98238 800
rect 98734 0 98790 800
rect 99286 0 99342 800
rect 99838 0 99894 800
rect 100390 0 100446 800
rect 100942 0 100998 800
rect 101494 0 101550 800
rect 102046 0 102102 800
rect 102598 0 102654 800
rect 103150 0 103206 800
rect 103702 0 103758 800
rect 104254 0 104310 800
rect 104806 0 104862 800
rect 105358 0 105414 800
rect 105910 0 105966 800
rect 106462 0 106518 800
rect 107014 0 107070 800
rect 107566 0 107622 800
rect 108118 0 108174 800
rect 108670 0 108726 800
rect 109222 0 109278 800
rect 109774 0 109830 800
rect 110326 0 110382 800
rect 110878 0 110934 800
rect 111430 0 111486 800
rect 111982 0 112038 800
rect 112534 0 112590 800
rect 113086 0 113142 800
rect 113638 0 113694 800
rect 114190 0 114246 800
rect 114742 0 114798 800
rect 115294 0 115350 800
rect 115846 0 115902 800
rect 116398 0 116454 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 118054 0 118110 800
rect 118606 0 118662 800
rect 119158 0 119214 800
rect 119710 0 119766 800
rect 120262 0 120318 800
rect 120814 0 120870 800
rect 121366 0 121422 800
rect 121918 0 121974 800
rect 122470 0 122526 800
rect 123022 0 123078 800
rect 123574 0 123630 800
rect 124126 0 124182 800
rect 124678 0 124734 800
rect 125230 0 125286 800
rect 125782 0 125838 800
rect 126334 0 126390 800
rect 126886 0 126942 800
rect 127438 0 127494 800
rect 127990 0 128046 800
rect 128542 0 128598 800
rect 129094 0 129150 800
rect 129646 0 129702 800
rect 130198 0 130254 800
rect 130750 0 130806 800
rect 131302 0 131358 800
rect 131854 0 131910 800
rect 132406 0 132462 800
rect 132958 0 133014 800
rect 133510 0 133566 800
rect 134062 0 134118 800
rect 134614 0 134670 800
rect 135166 0 135222 800
rect 135718 0 135774 800
rect 136270 0 136326 800
rect 136822 0 136878 800
rect 137374 0 137430 800
rect 137926 0 137982 800
rect 138478 0 138534 800
rect 139030 0 139086 800
rect 139582 0 139638 800
rect 140134 0 140190 800
rect 140686 0 140742 800
rect 141238 0 141294 800
rect 141790 0 141846 800
rect 142342 0 142398 800
rect 142894 0 142950 800
rect 143446 0 143502 800
rect 143998 0 144054 800
rect 144550 0 144606 800
rect 145102 0 145158 800
rect 145654 0 145710 800
rect 146206 0 146262 800
rect 146758 0 146814 800
rect 147310 0 147366 800
rect 147862 0 147918 800
rect 148414 0 148470 800
rect 148966 0 149022 800
rect 149518 0 149574 800
rect 150070 0 150126 800
rect 150622 0 150678 800
rect 151174 0 151230 800
rect 151726 0 151782 800
rect 152278 0 152334 800
rect 152830 0 152886 800
rect 153382 0 153438 800
rect 153934 0 153990 800
rect 154486 0 154542 800
rect 155038 0 155094 800
rect 155590 0 155646 800
rect 156142 0 156198 800
rect 156694 0 156750 800
rect 157246 0 157302 800
rect 157798 0 157854 800
rect 158350 0 158406 800
rect 158902 0 158958 800
rect 159454 0 159510 800
rect 160006 0 160062 800
rect 160558 0 160614 800
rect 161110 0 161166 800
rect 161662 0 161718 800
rect 162214 0 162270 800
rect 162766 0 162822 800
rect 163318 0 163374 800
rect 163870 0 163926 800
rect 164422 0 164478 800
rect 164974 0 165030 800
rect 165526 0 165582 800
rect 166078 0 166134 800
rect 166630 0 166686 800
rect 167182 0 167238 800
rect 167734 0 167790 800
rect 168286 0 168342 800
rect 168838 0 168894 800
rect 169390 0 169446 800
rect 169942 0 169998 800
rect 170494 0 170550 800
rect 171046 0 171102 800
rect 171598 0 171654 800
rect 172150 0 172206 800
rect 172702 0 172758 800
<< obsm2 >>
rect 3258 119144 4654 119354
rect 4822 119144 6218 119354
rect 6386 119144 7782 119354
rect 7950 119144 9346 119354
rect 9514 119144 10910 119354
rect 11078 119144 12474 119354
rect 12642 119144 14038 119354
rect 14206 119144 15602 119354
rect 15770 119144 17166 119354
rect 17334 119144 18730 119354
rect 18898 119144 20294 119354
rect 20462 119144 21858 119354
rect 22026 119144 23422 119354
rect 23590 119144 24986 119354
rect 25154 119144 26550 119354
rect 26718 119144 28114 119354
rect 28282 119144 29678 119354
rect 29846 119144 31242 119354
rect 31410 119144 32806 119354
rect 32974 119144 34370 119354
rect 34538 119144 35934 119354
rect 36102 119144 37498 119354
rect 37666 119144 39062 119354
rect 39230 119144 40626 119354
rect 40794 119144 42190 119354
rect 42358 119144 43754 119354
rect 43922 119144 45318 119354
rect 45486 119144 46882 119354
rect 47050 119144 48446 119354
rect 48614 119144 50010 119354
rect 50178 119144 51574 119354
rect 51742 119144 53138 119354
rect 53306 119144 54702 119354
rect 54870 119144 56266 119354
rect 56434 119144 57830 119354
rect 57998 119144 59394 119354
rect 59562 119144 60958 119354
rect 61126 119144 62522 119354
rect 62690 119144 64086 119354
rect 64254 119144 65650 119354
rect 65818 119144 67214 119354
rect 67382 119144 68778 119354
rect 68946 119144 70342 119354
rect 70510 119144 71906 119354
rect 72074 119144 73470 119354
rect 73638 119144 75034 119354
rect 75202 119144 76598 119354
rect 76766 119144 78162 119354
rect 78330 119144 79726 119354
rect 79894 119144 81290 119354
rect 81458 119144 82854 119354
rect 83022 119144 84418 119354
rect 84586 119144 85982 119354
rect 86150 119144 87546 119354
rect 87714 119144 89110 119354
rect 89278 119144 90674 119354
rect 90842 119144 92238 119354
rect 92406 119144 93802 119354
rect 93970 119144 95366 119354
rect 95534 119144 96930 119354
rect 97098 119144 98494 119354
rect 98662 119144 100058 119354
rect 100226 119144 101622 119354
rect 101790 119144 103186 119354
rect 103354 119144 104750 119354
rect 104918 119144 106314 119354
rect 106482 119144 107878 119354
rect 108046 119144 109442 119354
rect 109610 119144 111006 119354
rect 111174 119144 112570 119354
rect 112738 119144 114134 119354
rect 114302 119144 115698 119354
rect 115866 119144 117262 119354
rect 117430 119144 118826 119354
rect 118994 119144 120390 119354
rect 120558 119144 121954 119354
rect 122122 119144 123518 119354
rect 123686 119144 125082 119354
rect 125250 119144 126646 119354
rect 126814 119144 128210 119354
rect 128378 119144 129774 119354
rect 129942 119144 131338 119354
rect 131506 119144 132902 119354
rect 133070 119144 134466 119354
rect 134634 119144 136030 119354
rect 136198 119144 137594 119354
rect 137762 119144 139158 119354
rect 139326 119144 140722 119354
rect 140890 119144 142286 119354
rect 142454 119144 143850 119354
rect 144018 119144 145414 119354
rect 145582 119144 146978 119354
rect 147146 119144 148542 119354
rect 148710 119144 150106 119354
rect 150274 119144 151670 119354
rect 151838 119144 153234 119354
rect 153402 119144 154798 119354
rect 154966 119144 156362 119354
rect 156530 119144 157926 119354
rect 158094 119144 159490 119354
rect 159658 119144 161054 119354
rect 161222 119144 162618 119354
rect 162786 119144 164182 119354
rect 164350 119144 165746 119354
rect 165914 119144 167310 119354
rect 167478 119144 168874 119354
rect 169042 119144 170438 119354
rect 170606 119144 172002 119354
rect 172170 119144 173566 119354
rect 173734 119144 175130 119354
rect 175298 119144 176694 119354
rect 176862 119144 178258 119354
rect 3148 856 178368 119144
rect 3148 206 7046 856
rect 7214 206 7598 856
rect 7766 206 8150 856
rect 8318 206 8702 856
rect 8870 206 9254 856
rect 9422 206 9806 856
rect 9974 206 10358 856
rect 10526 206 10910 856
rect 11078 206 11462 856
rect 11630 206 12014 856
rect 12182 206 12566 856
rect 12734 206 13118 856
rect 13286 206 13670 856
rect 13838 206 14222 856
rect 14390 206 14774 856
rect 14942 206 15326 856
rect 15494 206 15878 856
rect 16046 206 16430 856
rect 16598 206 16982 856
rect 17150 206 17534 856
rect 17702 206 18086 856
rect 18254 206 18638 856
rect 18806 206 19190 856
rect 19358 206 19742 856
rect 19910 206 20294 856
rect 20462 206 20846 856
rect 21014 206 21398 856
rect 21566 206 21950 856
rect 22118 206 22502 856
rect 22670 206 23054 856
rect 23222 206 23606 856
rect 23774 206 24158 856
rect 24326 206 24710 856
rect 24878 206 25262 856
rect 25430 206 25814 856
rect 25982 206 26366 856
rect 26534 206 26918 856
rect 27086 206 27470 856
rect 27638 206 28022 856
rect 28190 206 28574 856
rect 28742 206 29126 856
rect 29294 206 29678 856
rect 29846 206 30230 856
rect 30398 206 30782 856
rect 30950 206 31334 856
rect 31502 206 31886 856
rect 32054 206 32438 856
rect 32606 206 32990 856
rect 33158 206 33542 856
rect 33710 206 34094 856
rect 34262 206 34646 856
rect 34814 206 35198 856
rect 35366 206 35750 856
rect 35918 206 36302 856
rect 36470 206 36854 856
rect 37022 206 37406 856
rect 37574 206 37958 856
rect 38126 206 38510 856
rect 38678 206 39062 856
rect 39230 206 39614 856
rect 39782 206 40166 856
rect 40334 206 40718 856
rect 40886 206 41270 856
rect 41438 206 41822 856
rect 41990 206 42374 856
rect 42542 206 42926 856
rect 43094 206 43478 856
rect 43646 206 44030 856
rect 44198 206 44582 856
rect 44750 206 45134 856
rect 45302 206 45686 856
rect 45854 206 46238 856
rect 46406 206 46790 856
rect 46958 206 47342 856
rect 47510 206 47894 856
rect 48062 206 48446 856
rect 48614 206 48998 856
rect 49166 206 49550 856
rect 49718 206 50102 856
rect 50270 206 50654 856
rect 50822 206 51206 856
rect 51374 206 51758 856
rect 51926 206 52310 856
rect 52478 206 52862 856
rect 53030 206 53414 856
rect 53582 206 53966 856
rect 54134 206 54518 856
rect 54686 206 55070 856
rect 55238 206 55622 856
rect 55790 206 56174 856
rect 56342 206 56726 856
rect 56894 206 57278 856
rect 57446 206 57830 856
rect 57998 206 58382 856
rect 58550 206 58934 856
rect 59102 206 59486 856
rect 59654 206 60038 856
rect 60206 206 60590 856
rect 60758 206 61142 856
rect 61310 206 61694 856
rect 61862 206 62246 856
rect 62414 206 62798 856
rect 62966 206 63350 856
rect 63518 206 63902 856
rect 64070 206 64454 856
rect 64622 206 65006 856
rect 65174 206 65558 856
rect 65726 206 66110 856
rect 66278 206 66662 856
rect 66830 206 67214 856
rect 67382 206 67766 856
rect 67934 206 68318 856
rect 68486 206 68870 856
rect 69038 206 69422 856
rect 69590 206 69974 856
rect 70142 206 70526 856
rect 70694 206 71078 856
rect 71246 206 71630 856
rect 71798 206 72182 856
rect 72350 206 72734 856
rect 72902 206 73286 856
rect 73454 206 73838 856
rect 74006 206 74390 856
rect 74558 206 74942 856
rect 75110 206 75494 856
rect 75662 206 76046 856
rect 76214 206 76598 856
rect 76766 206 77150 856
rect 77318 206 77702 856
rect 77870 206 78254 856
rect 78422 206 78806 856
rect 78974 206 79358 856
rect 79526 206 79910 856
rect 80078 206 80462 856
rect 80630 206 81014 856
rect 81182 206 81566 856
rect 81734 206 82118 856
rect 82286 206 82670 856
rect 82838 206 83222 856
rect 83390 206 83774 856
rect 83942 206 84326 856
rect 84494 206 84878 856
rect 85046 206 85430 856
rect 85598 206 85982 856
rect 86150 206 86534 856
rect 86702 206 87086 856
rect 87254 206 87638 856
rect 87806 206 88190 856
rect 88358 206 88742 856
rect 88910 206 89294 856
rect 89462 206 89846 856
rect 90014 206 90398 856
rect 90566 206 90950 856
rect 91118 206 91502 856
rect 91670 206 92054 856
rect 92222 206 92606 856
rect 92774 206 93158 856
rect 93326 206 93710 856
rect 93878 206 94262 856
rect 94430 206 94814 856
rect 94982 206 95366 856
rect 95534 206 95918 856
rect 96086 206 96470 856
rect 96638 206 97022 856
rect 97190 206 97574 856
rect 97742 206 98126 856
rect 98294 206 98678 856
rect 98846 206 99230 856
rect 99398 206 99782 856
rect 99950 206 100334 856
rect 100502 206 100886 856
rect 101054 206 101438 856
rect 101606 206 101990 856
rect 102158 206 102542 856
rect 102710 206 103094 856
rect 103262 206 103646 856
rect 103814 206 104198 856
rect 104366 206 104750 856
rect 104918 206 105302 856
rect 105470 206 105854 856
rect 106022 206 106406 856
rect 106574 206 106958 856
rect 107126 206 107510 856
rect 107678 206 108062 856
rect 108230 206 108614 856
rect 108782 206 109166 856
rect 109334 206 109718 856
rect 109886 206 110270 856
rect 110438 206 110822 856
rect 110990 206 111374 856
rect 111542 206 111926 856
rect 112094 206 112478 856
rect 112646 206 113030 856
rect 113198 206 113582 856
rect 113750 206 114134 856
rect 114302 206 114686 856
rect 114854 206 115238 856
rect 115406 206 115790 856
rect 115958 206 116342 856
rect 116510 206 116894 856
rect 117062 206 117446 856
rect 117614 206 117998 856
rect 118166 206 118550 856
rect 118718 206 119102 856
rect 119270 206 119654 856
rect 119822 206 120206 856
rect 120374 206 120758 856
rect 120926 206 121310 856
rect 121478 206 121862 856
rect 122030 206 122414 856
rect 122582 206 122966 856
rect 123134 206 123518 856
rect 123686 206 124070 856
rect 124238 206 124622 856
rect 124790 206 125174 856
rect 125342 206 125726 856
rect 125894 206 126278 856
rect 126446 206 126830 856
rect 126998 206 127382 856
rect 127550 206 127934 856
rect 128102 206 128486 856
rect 128654 206 129038 856
rect 129206 206 129590 856
rect 129758 206 130142 856
rect 130310 206 130694 856
rect 130862 206 131246 856
rect 131414 206 131798 856
rect 131966 206 132350 856
rect 132518 206 132902 856
rect 133070 206 133454 856
rect 133622 206 134006 856
rect 134174 206 134558 856
rect 134726 206 135110 856
rect 135278 206 135662 856
rect 135830 206 136214 856
rect 136382 206 136766 856
rect 136934 206 137318 856
rect 137486 206 137870 856
rect 138038 206 138422 856
rect 138590 206 138974 856
rect 139142 206 139526 856
rect 139694 206 140078 856
rect 140246 206 140630 856
rect 140798 206 141182 856
rect 141350 206 141734 856
rect 141902 206 142286 856
rect 142454 206 142838 856
rect 143006 206 143390 856
rect 143558 206 143942 856
rect 144110 206 144494 856
rect 144662 206 145046 856
rect 145214 206 145598 856
rect 145766 206 146150 856
rect 146318 206 146702 856
rect 146870 206 147254 856
rect 147422 206 147806 856
rect 147974 206 148358 856
rect 148526 206 148910 856
rect 149078 206 149462 856
rect 149630 206 150014 856
rect 150182 206 150566 856
rect 150734 206 151118 856
rect 151286 206 151670 856
rect 151838 206 152222 856
rect 152390 206 152774 856
rect 152942 206 153326 856
rect 153494 206 153878 856
rect 154046 206 154430 856
rect 154598 206 154982 856
rect 155150 206 155534 856
rect 155702 206 156086 856
rect 156254 206 156638 856
rect 156806 206 157190 856
rect 157358 206 157742 856
rect 157910 206 158294 856
rect 158462 206 158846 856
rect 159014 206 159398 856
rect 159566 206 159950 856
rect 160118 206 160502 856
rect 160670 206 161054 856
rect 161222 206 161606 856
rect 161774 206 162158 856
rect 162326 206 162710 856
rect 162878 206 163262 856
rect 163430 206 163814 856
rect 163982 206 164366 856
rect 164534 206 164918 856
rect 165086 206 165470 856
rect 165638 206 166022 856
rect 166190 206 166574 856
rect 166742 206 167126 856
rect 167294 206 167678 856
rect 167846 206 168230 856
rect 168398 206 168782 856
rect 168950 206 169334 856
rect 169502 206 169886 856
rect 170054 206 170438 856
rect 170606 206 170990 856
rect 171158 206 171542 856
rect 171710 206 172094 856
rect 172262 206 172646 856
rect 172814 206 178368 856
<< obsm3 >>
rect 4210 443 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 77339 2048 80928 8397
rect 81408 2048 96288 8397
rect 96768 2048 111648 8397
rect 112128 2048 126533 8397
rect 77339 443 126533 2048
<< labels >>
rlabel metal2 s 1582 119200 1638 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 48502 119200 48558 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 53194 119200 53250 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57886 119200 57942 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 62578 119200 62634 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 67270 119200 67326 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71962 119200 72018 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 76654 119200 76710 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81346 119200 81402 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86038 119200 86094 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 90730 119200 90786 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6274 119200 6330 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95422 119200 95478 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100114 119200 100170 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104806 119200 104862 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 109498 119200 109554 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114190 119200 114246 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118882 119200 118938 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 123574 119200 123630 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 128266 119200 128322 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 132958 119200 133014 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 137650 119200 137706 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10966 119200 11022 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 142342 119200 142398 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 147034 119200 147090 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 151726 119200 151782 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 156418 119200 156474 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 161110 119200 161166 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 165802 119200 165858 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 170494 119200 170550 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 175186 119200 175242 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 15658 119200 15714 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 20350 119200 20406 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 25042 119200 25098 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29734 119200 29790 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 34426 119200 34482 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 39118 119200 39174 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3146 119200 3202 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 50066 119200 50122 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 54758 119200 54814 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 59450 119200 59506 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 64142 119200 64198 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68834 119200 68890 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 73526 119200 73582 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 78218 119200 78274 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82910 119200 82966 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 87602 119200 87658 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92294 119200 92350 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7838 119200 7894 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 96986 119200 97042 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 101678 119200 101734 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 111062 119200 111118 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 115754 119200 115810 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 120446 119200 120502 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 125138 119200 125194 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 129830 119200 129886 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 134522 119200 134578 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 139214 119200 139270 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12530 119200 12586 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 143906 119200 143962 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 148598 119200 148654 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 153290 119200 153346 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 157982 119200 158038 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 162674 119200 162730 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 167366 119200 167422 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 172058 119200 172114 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 176750 119200 176806 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 17222 119200 17278 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21914 119200 21970 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 26606 119200 26662 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 31298 119200 31354 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35990 119200 36046 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 40682 119200 40738 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 45374 119200 45430 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4710 119200 4766 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 51630 119200 51686 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 56322 119200 56378 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 61014 119200 61070 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 65706 119200 65762 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 70398 119200 70454 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 79782 119200 79838 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 84474 119200 84530 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 89166 119200 89222 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93858 119200 93914 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9402 119200 9458 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 98550 119200 98606 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 103242 119200 103298 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 107934 119200 107990 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 112626 119200 112682 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 117318 119200 117374 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 122010 119200 122066 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 126702 119200 126758 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 131394 119200 131450 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 136086 119200 136142 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 140778 119200 140834 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14094 119200 14150 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 145470 119200 145526 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 150162 119200 150218 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 154854 119200 154910 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 159546 119200 159602 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 164238 119200 164294 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 168930 119200 168986 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 173622 119200 173678 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 178314 119200 178370 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18786 119200 18842 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 23478 119200 23534 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 28170 119200 28226 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32862 119200 32918 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37554 119200 37610 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 42246 119200 42302 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46938 119200 46994 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 172150 0 172206 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[32]
port 143 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[35]
port 146 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[38]
port 149 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[39]
port 150 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[3]
port 151 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[40]
port 152 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[41]
port 153 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[48]
port 160 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[4]
port 162 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[50]
port 163 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[51]
port 164 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[52]
port 165 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[54]
port 167 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[59]
port 172 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_data_in[60]
port 174 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[6]
port 178 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[8]
port 180 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_out[0]
port 182 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[10]
port 183 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[11]
port 184 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[15]
port 188 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[17]
port 190 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[18]
port 191 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[1]
port 193 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[20]
port 194 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[21]
port 195 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[23]
port 197 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 la_data_out[25]
port 199 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[26]
port 200 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 la_data_out[27]
port 201 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[29]
port 203 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[31]
port 206 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[32]
port 207 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_out[33]
port 208 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 la_data_out[34]
port 209 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_data_out[35]
port 210 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 la_data_out[36]
port 211 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[37]
port 212 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[38]
port 213 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 la_data_out[42]
port 218 nsew signal output
rlabel metal2 s 137374 0 137430 800 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 la_data_out[47]
port 223 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 la_data_out[49]
port 225 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[51]
port 228 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[52]
port 229 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[53]
port 230 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[54]
port 231 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[55]
port 232 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 160558 0 160614 800 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[59]
port 236 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[5]
port 237 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 167182 0 167238 800 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 168838 0 168894 800 6 la_data_out[62]
port 240 nsew signal output
rlabel metal2 s 170494 0 170550 800 6 la_data_out[63]
port 241 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[6]
port 242 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[7]
port 243 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[12]
port 249 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[14]
port 251 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[16]
port 253 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[1]
port 257 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[21]
port 259 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[23]
port 261 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[24]
port 262 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_oenb[26]
port 264 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[27]
port 265 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[28]
port 266 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[34]
port 273 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_oenb[35]
port 274 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oenb[36]
port 275 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[38]
port 277 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[40]
port 280 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[43]
port 283 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_oenb[44]
port 284 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[45]
port 285 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oenb[49]
port 289 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[50]
port 291 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_oenb[53]
port 294 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_oenb[56]
port 297 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[58]
port 299 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[59]
port 300 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[5]
port 301 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_oenb[62]
port 304 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oenb[6]
port 306 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[8]
port 308 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 310 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 310 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 310 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 310 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 310 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 310 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 311 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 311 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 311 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 311 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 311 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 311 nsew ground bidirectional
rlabel metal2 s 7102 0 7158 800 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wb_rst_i
port 313 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_stb_i
port 416 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7897226
string GDS_FILE /home/mpotereau/DigitalFlowTest/gf_spi_test/openlane/user_proj_example/runs/23_01_09_10_45/results/signoff/user_proj_example.magic.gds
string GDS_START 350044
<< end >>

