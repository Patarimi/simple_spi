magic
tech sky130A
magscale 1 2
timestamp 1673535535
<< viali >>
rect 1777 15657 1811 15691
rect 4353 15657 4387 15691
rect 7757 15657 7791 15691
rect 10701 15657 10735 15691
rect 16221 15657 16255 15691
rect 1961 15453 1995 15487
rect 2421 15453 2455 15487
rect 3249 15453 3283 15487
rect 4537 15453 4571 15487
rect 5733 15453 5767 15487
rect 6009 15453 6043 15487
rect 6745 15453 6779 15487
rect 7573 15453 7607 15487
rect 10517 15453 10551 15487
rect 16037 15453 16071 15487
rect 2513 15385 2547 15419
rect 3157 15317 3191 15351
rect 4997 15317 5031 15351
rect 6561 15317 6595 15351
rect 1593 15113 1627 15147
rect 8217 15113 8251 15147
rect 2329 14977 2363 15011
rect 2605 14977 2639 15011
rect 5549 14977 5583 15011
rect 5641 14977 5675 15011
rect 5825 14977 5859 15011
rect 7481 14977 7515 15011
rect 3065 14909 3099 14943
rect 3341 14909 3375 14943
rect 5089 14909 5123 14943
rect 6009 14909 6043 14943
rect 7205 14909 7239 14943
rect 6561 14841 6595 14875
rect 7297 14569 7331 14603
rect 4261 14433 4295 14467
rect 3433 14365 3467 14399
rect 3985 14365 4019 14399
rect 6285 14365 6319 14399
rect 6561 14365 6595 14399
rect 7757 14365 7791 14399
rect 8033 14365 8067 14399
rect 8217 14297 8251 14331
rect 2145 14229 2179 14263
rect 5733 14229 5767 14263
rect 7849 14229 7883 14263
rect 1860 14025 1894 14059
rect 6009 13957 6043 13991
rect 1593 13889 1627 13923
rect 2237 13889 2271 13923
rect 5549 13889 5583 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 7021 13889 7055 13923
rect 7113 13889 7147 13923
rect 7205 13889 7239 13923
rect 3157 13821 3191 13855
rect 3433 13821 3467 13855
rect 6837 13821 6871 13855
rect 1869 13685 1903 13719
rect 4905 13685 4939 13719
rect 6285 13481 6319 13515
rect 7297 13481 7331 13515
rect 7481 13481 7515 13515
rect 1593 13345 1627 13379
rect 1869 13345 1903 13379
rect 3341 13345 3375 13379
rect 5733 13345 5767 13379
rect 7205 13345 7239 13379
rect 3985 13277 4019 13311
rect 6193 13277 6227 13311
rect 6929 13277 6963 13311
rect 4261 13209 4295 13243
rect 2053 12937 2087 12971
rect 3893 12937 3927 12971
rect 6561 12937 6595 12971
rect 2605 12869 2639 12903
rect 1961 12801 1995 12835
rect 5089 12801 5123 12835
rect 5181 12801 5215 12835
rect 5365 12801 5399 12835
rect 6745 12801 6779 12835
rect 7113 12801 7147 12835
rect 5273 12733 5307 12767
rect 5549 12597 5583 12631
rect 7021 12597 7055 12631
rect 4629 12393 4663 12427
rect 1593 12257 1627 12291
rect 5549 12257 5583 12291
rect 5917 12257 5951 12291
rect 3341 12189 3375 12223
rect 4169 12189 4203 12223
rect 4813 12189 4847 12223
rect 5457 12189 5491 12223
rect 6377 12189 6411 12223
rect 6745 12189 6779 12223
rect 8309 12189 8343 12223
rect 6561 12121 6595 12155
rect 3985 12053 4019 12087
rect 5273 12053 5307 12087
rect 8493 12053 8527 12087
rect 3433 11849 3467 11883
rect 5089 11849 5123 11883
rect 5273 11849 5307 11883
rect 2329 11713 2363 11747
rect 3617 11713 3651 11747
rect 3893 11713 3927 11747
rect 4077 11713 4111 11747
rect 5270 11713 5304 11747
rect 6561 11713 6595 11747
rect 8585 11713 8619 11747
rect 8861 11713 8895 11747
rect 2605 11645 2639 11679
rect 5733 11645 5767 11679
rect 1593 11509 1627 11543
rect 5641 11509 5675 11543
rect 6745 11509 6779 11543
rect 9597 11509 9631 11543
rect 2789 11305 2823 11339
rect 4067 11305 4101 11339
rect 1869 11237 1903 11271
rect 3249 11237 3283 11271
rect 5549 11237 5583 11271
rect 5917 11237 5951 11271
rect 6009 11169 6043 11203
rect 1685 11101 1719 11135
rect 2605 11101 2639 11135
rect 3433 11101 3467 11135
rect 4813 11101 4847 11135
rect 5089 11101 5123 11135
rect 5733 11101 5767 11135
rect 2789 10761 2823 10795
rect 4169 10761 4203 10795
rect 5549 10761 5583 10795
rect 6561 10761 6595 10795
rect 1961 10693 1995 10727
rect 2145 10625 2179 10659
rect 2329 10625 2363 10659
rect 3709 10625 3743 10659
rect 5365 10625 5399 10659
rect 6745 10625 6779 10659
rect 6837 10625 6871 10659
rect 6929 10625 6963 10659
rect 3985 10421 4019 10455
rect 1777 10217 1811 10251
rect 4353 10217 4387 10251
rect 4537 10217 4571 10251
rect 7113 10217 7147 10251
rect 3985 10149 4019 10183
rect 7389 10081 7423 10115
rect 1869 10013 1903 10047
rect 7481 10013 7515 10047
rect 4353 9945 4387 9979
rect 2237 9537 2271 9571
rect 4077 9537 4111 9571
rect 3801 9469 3835 9503
rect 2421 9401 2455 9435
rect 3525 9333 3559 9367
rect 3709 9333 3743 9367
rect 2053 9129 2087 9163
rect 1869 8925 1903 8959
rect 1593 6749 1627 6783
rect 2237 6749 2271 6783
rect 1777 6613 1811 6647
rect 1593 2397 1627 2431
rect 1777 2261 1811 2295
<< metal1 >>
rect 1104 15802 16836 15824
rect 1104 15750 2916 15802
rect 2968 15750 2980 15802
rect 3032 15750 3044 15802
rect 3096 15750 3108 15802
rect 3160 15750 3172 15802
rect 3224 15750 6849 15802
rect 6901 15750 6913 15802
rect 6965 15750 6977 15802
rect 7029 15750 7041 15802
rect 7093 15750 7105 15802
rect 7157 15750 10782 15802
rect 10834 15750 10846 15802
rect 10898 15750 10910 15802
rect 10962 15750 10974 15802
rect 11026 15750 11038 15802
rect 11090 15750 14715 15802
rect 14767 15750 14779 15802
rect 14831 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 16836 15802
rect 1104 15728 16836 15750
rect 1578 15648 1584 15700
rect 1636 15688 1642 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1636 15660 1777 15688
rect 1636 15648 1642 15660
rect 1765 15657 1777 15660
rect 1811 15657 1823 15691
rect 1765 15651 1823 15657
rect 4341 15691 4399 15697
rect 4341 15657 4353 15691
rect 4387 15688 4399 15691
rect 4522 15688 4528 15700
rect 4387 15660 4528 15688
rect 4387 15657 4399 15660
rect 4341 15651 4399 15657
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 7745 15691 7803 15697
rect 7745 15688 7757 15691
rect 7524 15660 7757 15688
rect 7524 15648 7530 15660
rect 7745 15657 7757 15660
rect 7791 15657 7803 15691
rect 10686 15688 10692 15700
rect 10647 15660 10692 15688
rect 7745 15651 7803 15657
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 16206 15688 16212 15700
rect 16167 15660 16212 15688
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 3786 15620 3792 15632
rect 1964 15592 3792 15620
rect 1964 15493 1992 15592
rect 3786 15580 3792 15592
rect 3844 15580 3850 15632
rect 2038 15512 2044 15564
rect 2096 15552 2102 15564
rect 2096 15524 5396 15552
rect 2096 15512 2102 15524
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15453 2007 15487
rect 2406 15484 2412 15496
rect 2367 15456 2412 15484
rect 1949 15447 2007 15453
rect 2406 15444 2412 15456
rect 2464 15484 2470 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 2464 15456 3249 15484
rect 2464 15444 2470 15456
rect 3237 15453 3249 15456
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 4571 15456 5028 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 2501 15419 2559 15425
rect 2501 15385 2513 15419
rect 2547 15416 2559 15419
rect 3694 15416 3700 15428
rect 2547 15388 3700 15416
rect 2547 15385 2559 15388
rect 2501 15379 2559 15385
rect 3694 15376 3700 15388
rect 3752 15376 3758 15428
rect 3145 15351 3203 15357
rect 3145 15317 3157 15351
rect 3191 15348 3203 15351
rect 3234 15348 3240 15360
rect 3191 15320 3240 15348
rect 3191 15317 3203 15320
rect 3145 15311 3203 15317
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 5000 15357 5028 15456
rect 5368 15416 5396 15524
rect 5718 15484 5724 15496
rect 5679 15456 5724 15484
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 5994 15484 6000 15496
rect 5955 15456 6000 15484
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 7558 15484 7564 15496
rect 7519 15456 7564 15484
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 8352 15456 10517 15484
rect 8352 15444 8358 15456
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 16025 15487 16083 15493
rect 16025 15453 16037 15487
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 16040 15416 16068 15447
rect 5368 15388 16068 15416
rect 4985 15351 5043 15357
rect 4985 15317 4997 15351
rect 5031 15317 5043 15351
rect 6546 15348 6552 15360
rect 6507 15320 6552 15348
rect 4985 15311 5043 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 1104 15258 16995 15280
rect 1104 15206 4882 15258
rect 4934 15206 4946 15258
rect 4998 15206 5010 15258
rect 5062 15206 5074 15258
rect 5126 15206 5138 15258
rect 5190 15206 8815 15258
rect 8867 15206 8879 15258
rect 8931 15206 8943 15258
rect 8995 15206 9007 15258
rect 9059 15206 9071 15258
rect 9123 15206 12748 15258
rect 12800 15206 12812 15258
rect 12864 15206 12876 15258
rect 12928 15206 12940 15258
rect 12992 15206 13004 15258
rect 13056 15206 16681 15258
rect 16733 15206 16745 15258
rect 16797 15206 16809 15258
rect 16861 15206 16873 15258
rect 16925 15206 16937 15258
rect 16989 15206 16995 15258
rect 1104 15184 16995 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 2038 15144 2044 15156
rect 1627 15116 2044 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 6546 15144 6552 15156
rect 2332 15116 6552 15144
rect 2332 15017 2360 15116
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8294 15144 8300 15156
rect 8251 15116 8300 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 3602 15076 3608 15088
rect 2608 15048 3608 15076
rect 2608 15017 2636 15048
rect 3602 15036 3608 15048
rect 3660 15036 3666 15088
rect 6270 15076 6276 15088
rect 4554 15048 6276 15076
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 5442 14968 5448 15020
rect 5500 15008 5506 15020
rect 5537 15011 5595 15017
rect 5537 15008 5549 15011
rect 5500 14980 5549 15008
rect 5500 14968 5506 14980
rect 5537 14977 5549 14980
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 5684 14980 5729 15008
rect 5684 14968 5690 14980
rect 5810 14968 5816 15020
rect 5868 15008 5874 15020
rect 5868 14980 5913 15008
rect 5868 14968 5874 14980
rect 6546 14968 6552 15020
rect 6604 15008 6610 15020
rect 7469 15011 7527 15017
rect 7469 15008 7481 15011
rect 6604 14980 7481 15008
rect 6604 14968 6610 14980
rect 7469 14977 7481 14980
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 2682 14900 2688 14952
rect 2740 14940 2746 14952
rect 3053 14943 3111 14949
rect 3053 14940 3065 14943
rect 2740 14912 3065 14940
rect 2740 14900 2746 14912
rect 3053 14909 3065 14912
rect 3099 14909 3111 14943
rect 3326 14940 3332 14952
rect 3287 14912 3332 14940
rect 3053 14903 3111 14909
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5828 14940 5856 14968
rect 5123 14912 5856 14940
rect 5997 14943 6055 14949
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5997 14909 6009 14943
rect 6043 14940 6055 14943
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6043 14912 7205 14940
rect 6043 14909 6055 14912
rect 5997 14903 6055 14909
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 6549 14875 6607 14881
rect 6549 14872 6561 14875
rect 4356 14844 6561 14872
rect 2774 14764 2780 14816
rect 2832 14804 2838 14816
rect 4356 14804 4384 14844
rect 6549 14841 6561 14844
rect 6595 14841 6607 14875
rect 6549 14835 6607 14841
rect 2832 14776 4384 14804
rect 2832 14764 2838 14776
rect 1104 14714 16836 14736
rect 1104 14662 2916 14714
rect 2968 14662 2980 14714
rect 3032 14662 3044 14714
rect 3096 14662 3108 14714
rect 3160 14662 3172 14714
rect 3224 14662 6849 14714
rect 6901 14662 6913 14714
rect 6965 14662 6977 14714
rect 7029 14662 7041 14714
rect 7093 14662 7105 14714
rect 7157 14662 10782 14714
rect 10834 14662 10846 14714
rect 10898 14662 10910 14714
rect 10962 14662 10974 14714
rect 11026 14662 11038 14714
rect 11090 14662 14715 14714
rect 14767 14662 14779 14714
rect 14831 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 16836 14714
rect 1104 14640 16836 14662
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 6822 14600 6828 14612
rect 5868 14572 6828 14600
rect 5868 14560 5874 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 7558 14600 7564 14612
rect 7331 14572 7564 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 6840 14532 6868 14560
rect 6840 14504 8064 14532
rect 4249 14467 4307 14473
rect 4249 14433 4261 14467
rect 4295 14464 4307 14467
rect 5810 14464 5816 14476
rect 4295 14436 5816 14464
rect 4295 14433 4307 14436
rect 4249 14427 4307 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 2774 14356 2780 14408
rect 2832 14396 2838 14408
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 2832 14368 3433 14396
rect 2832 14356 2838 14368
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3936 14368 3985 14396
rect 3936 14356 3942 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 6546 14396 6552 14408
rect 6507 14368 6552 14396
rect 6273 14359 6331 14365
rect 6288 14328 6316 14359
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 7742 14396 7748 14408
rect 7703 14368 7748 14396
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 8036 14405 8064 14504
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8205 14331 8263 14337
rect 8205 14328 8217 14331
rect 4356 14300 4738 14328
rect 6288 14300 8217 14328
rect 2130 14260 2136 14272
rect 2091 14232 2136 14260
rect 2130 14220 2136 14232
rect 2188 14220 2194 14272
rect 3694 14220 3700 14272
rect 3752 14260 3758 14272
rect 4356 14260 4384 14300
rect 8205 14297 8217 14300
rect 8251 14297 8263 14331
rect 8205 14291 8263 14297
rect 3752 14232 4384 14260
rect 5721 14263 5779 14269
rect 3752 14220 3758 14232
rect 5721 14229 5733 14263
rect 5767 14260 5779 14263
rect 6638 14260 6644 14272
rect 5767 14232 6644 14260
rect 5767 14229 5779 14232
rect 5721 14223 5779 14229
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 7834 14260 7840 14272
rect 7795 14232 7840 14260
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 1104 14170 16995 14192
rect 1104 14118 4882 14170
rect 4934 14118 4946 14170
rect 4998 14118 5010 14170
rect 5062 14118 5074 14170
rect 5126 14118 5138 14170
rect 5190 14118 8815 14170
rect 8867 14118 8879 14170
rect 8931 14118 8943 14170
rect 8995 14118 9007 14170
rect 9059 14118 9071 14170
rect 9123 14118 12748 14170
rect 12800 14118 12812 14170
rect 12864 14118 12876 14170
rect 12928 14118 12940 14170
rect 12992 14118 13004 14170
rect 13056 14118 16681 14170
rect 16733 14118 16745 14170
rect 16797 14118 16809 14170
rect 16861 14118 16873 14170
rect 16925 14118 16937 14170
rect 16989 14118 16995 14170
rect 1104 14096 16995 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 1848 14059 1906 14065
rect 1848 14056 1860 14059
rect 1636 14028 1860 14056
rect 1636 14016 1642 14028
rect 1848 14025 1860 14028
rect 1894 14056 1906 14059
rect 2682 14056 2688 14068
rect 1894 14028 2688 14056
rect 1894 14025 1906 14028
rect 1848 14019 1906 14025
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 6730 14056 6736 14068
rect 3804 14028 6736 14056
rect 3804 13988 3832 14028
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 1596 13960 3832 13988
rect 1596 13929 1624 13960
rect 4154 13948 4160 14000
rect 4212 13948 4218 14000
rect 5718 13948 5724 14000
rect 5776 13988 5782 14000
rect 5994 13988 6000 14000
rect 5776 13960 5856 13988
rect 5955 13960 6000 13988
rect 5776 13948 5782 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 1581 13883 1639 13889
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 5534 13920 5540 13932
rect 5495 13892 5540 13920
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 5828 13929 5856 13960
rect 5994 13948 6000 13960
rect 6052 13948 6058 14000
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 6696 13960 7144 13988
rect 6696 13948 6702 13960
rect 7116 13929 7144 13960
rect 5813 13923 5871 13929
rect 5684 13892 5729 13920
rect 5684 13880 5690 13892
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 5813 13883 5871 13889
rect 5920 13892 7021 13920
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 3418 13852 3424 13864
rect 3191 13824 3280 13852
rect 3379 13824 3424 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 1857 13719 1915 13725
rect 1857 13685 1869 13719
rect 1903 13716 1915 13719
rect 2222 13716 2228 13728
rect 1903 13688 2228 13716
rect 1903 13685 1915 13688
rect 1857 13679 1915 13685
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 3252 13716 3280 13824
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 5920 13784 5948 13892
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 5276 13756 5948 13784
rect 6012 13824 6837 13852
rect 5276 13728 5304 13756
rect 3878 13716 3884 13728
rect 3252 13688 3884 13716
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 4893 13719 4951 13725
rect 4893 13685 4905 13719
rect 4939 13716 4951 13719
rect 5258 13716 5264 13728
rect 4939 13688 5264 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 5442 13676 5448 13728
rect 5500 13716 5506 13728
rect 6012 13716 6040 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 7024 13852 7052 13883
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7248 13892 7293 13920
rect 7248 13880 7254 13892
rect 7282 13852 7288 13864
rect 7024 13824 7288 13852
rect 6825 13815 6883 13821
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 5500 13688 6040 13716
rect 5500 13676 5506 13688
rect 1104 13626 16836 13648
rect 1104 13574 2916 13626
rect 2968 13574 2980 13626
rect 3032 13574 3044 13626
rect 3096 13574 3108 13626
rect 3160 13574 3172 13626
rect 3224 13574 6849 13626
rect 6901 13574 6913 13626
rect 6965 13574 6977 13626
rect 7029 13574 7041 13626
rect 7093 13574 7105 13626
rect 7157 13574 10782 13626
rect 10834 13574 10846 13626
rect 10898 13574 10910 13626
rect 10962 13574 10974 13626
rect 11026 13574 11038 13626
rect 11090 13574 14715 13626
rect 14767 13574 14779 13626
rect 14831 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 16836 13626
rect 1104 13552 16836 13574
rect 4430 13512 4436 13524
rect 3252 13484 4436 13512
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13376 1915 13379
rect 3252 13376 3280 13484
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 6270 13512 6276 13524
rect 6231 13484 6276 13512
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 7282 13512 7288 13524
rect 7243 13484 7288 13512
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7469 13515 7527 13521
rect 7469 13481 7481 13515
rect 7515 13512 7527 13515
rect 7742 13512 7748 13524
rect 7515 13484 7748 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 1903 13348 3280 13376
rect 3329 13379 3387 13385
rect 1903 13345 1915 13348
rect 1857 13339 1915 13345
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 4614 13376 4620 13388
rect 3375 13348 4620 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 5718 13376 5724 13388
rect 5631 13348 5724 13376
rect 5718 13336 5724 13348
rect 5776 13376 5782 13388
rect 7190 13376 7196 13388
rect 5776 13348 7196 13376
rect 5776 13336 5782 13348
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3936 13280 3985 13308
rect 3936 13268 3942 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 6178 13308 6184 13320
rect 6139 13280 6184 13308
rect 3973 13271 4031 13277
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6546 13308 6552 13320
rect 6328 13280 6552 13308
rect 6328 13268 6334 13280
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6696 13280 6929 13308
rect 6696 13268 6702 13280
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 3234 13240 3240 13252
rect 3082 13212 3240 13240
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 4246 13240 4252 13252
rect 4207 13212 4252 13240
rect 4246 13200 4252 13212
rect 4304 13200 4310 13252
rect 4356 13212 4738 13240
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 4356 13172 4384 13212
rect 3752 13144 4384 13172
rect 3752 13132 3758 13144
rect 1104 13082 16995 13104
rect 1104 13030 4882 13082
rect 4934 13030 4946 13082
rect 4998 13030 5010 13082
rect 5062 13030 5074 13082
rect 5126 13030 5138 13082
rect 5190 13030 8815 13082
rect 8867 13030 8879 13082
rect 8931 13030 8943 13082
rect 8995 13030 9007 13082
rect 9059 13030 9071 13082
rect 9123 13030 12748 13082
rect 12800 13030 12812 13082
rect 12864 13030 12876 13082
rect 12928 13030 12940 13082
rect 12992 13030 13004 13082
rect 13056 13030 16681 13082
rect 16733 13030 16745 13082
rect 16797 13030 16809 13082
rect 16861 13030 16873 13082
rect 16925 13030 16937 13082
rect 16989 13030 16995 13082
rect 1104 13008 16995 13030
rect 2041 12971 2099 12977
rect 2041 12937 2053 12971
rect 2087 12968 2099 12971
rect 3694 12968 3700 12980
rect 2087 12940 3700 12968
rect 2087 12937 2099 12940
rect 2041 12931 2099 12937
rect 3694 12928 3700 12940
rect 3752 12928 3758 12980
rect 3878 12968 3884 12980
rect 3839 12940 3884 12968
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 5592 12940 6561 12968
rect 5592 12928 5598 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 2130 12860 2136 12912
rect 2188 12900 2194 12912
rect 2590 12900 2596 12912
rect 2188 12872 2596 12900
rect 2188 12860 2194 12872
rect 2590 12860 2596 12872
rect 2648 12860 2654 12912
rect 6178 12900 6184 12912
rect 2746 12872 6184 12900
rect 1854 12792 1860 12844
rect 1912 12832 1918 12844
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1912 12804 1961 12832
rect 1912 12792 1918 12804
rect 1949 12801 1961 12804
rect 1995 12832 2007 12835
rect 2406 12832 2412 12844
rect 1995 12804 2412 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2406 12792 2412 12804
rect 2464 12832 2470 12844
rect 2746 12832 2774 12872
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 2464 12804 2774 12832
rect 2464 12792 2470 12804
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 4798 12832 4804 12844
rect 4672 12804 4804 12832
rect 4672 12792 4678 12804
rect 4798 12792 4804 12804
rect 4856 12832 4862 12844
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4856 12804 5089 12832
rect 4856 12792 4862 12804
rect 5077 12801 5089 12804
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5353 12835 5411 12841
rect 5224 12804 5269 12832
rect 5224 12792 5230 12804
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5626 12832 5632 12844
rect 5399 12804 5632 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5626 12792 5632 12804
rect 5684 12832 5690 12844
rect 6638 12832 6644 12844
rect 5684 12804 6644 12832
rect 5684 12792 5690 12804
rect 6638 12792 6644 12804
rect 6696 12832 6702 12844
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 6696 12804 6745 12832
rect 6696 12792 6702 12804
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 7282 12832 7288 12844
rect 7147 12804 7288 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12764 5319 12767
rect 5718 12764 5724 12776
rect 5307 12736 5724 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 6748 12764 6776 12795
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7466 12764 7472 12776
rect 6748 12736 7472 12764
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 5537 12631 5595 12637
rect 5537 12597 5549 12631
rect 5583 12628 5595 12631
rect 6362 12628 6368 12640
rect 5583 12600 6368 12628
rect 5583 12597 5595 12600
rect 5537 12591 5595 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7190 12628 7196 12640
rect 7055 12600 7196 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 1104 12538 16836 12560
rect 1104 12486 2916 12538
rect 2968 12486 2980 12538
rect 3032 12486 3044 12538
rect 3096 12486 3108 12538
rect 3160 12486 3172 12538
rect 3224 12486 6849 12538
rect 6901 12486 6913 12538
rect 6965 12486 6977 12538
rect 7029 12486 7041 12538
rect 7093 12486 7105 12538
rect 7157 12486 10782 12538
rect 10834 12486 10846 12538
rect 10898 12486 10910 12538
rect 10962 12486 10974 12538
rect 11026 12486 11038 12538
rect 11090 12486 14715 12538
rect 14767 12486 14779 12538
rect 14831 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 16836 12538
rect 1104 12464 16836 12486
rect 4614 12424 4620 12436
rect 4575 12396 4620 12424
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 1578 12288 1584 12300
rect 1539 12260 1584 12288
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 5537 12291 5595 12297
rect 5537 12257 5549 12291
rect 5583 12288 5595 12291
rect 5626 12288 5632 12300
rect 5583 12260 5632 12288
rect 5583 12257 5595 12260
rect 5537 12251 5595 12257
rect 5626 12248 5632 12260
rect 5684 12248 5690 12300
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5776 12260 5917 12288
rect 5776 12248 5782 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 2590 12180 2596 12232
rect 2648 12220 2654 12232
rect 3329 12223 3387 12229
rect 3329 12220 3341 12223
rect 2648 12192 3341 12220
rect 2648 12180 2654 12192
rect 3329 12189 3341 12192
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 4120 12192 4169 12220
rect 4120 12180 4126 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4798 12220 4804 12232
rect 4759 12192 4804 12220
rect 4157 12183 4215 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5350 12180 5356 12232
rect 5408 12220 5414 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5408 12192 5457 12220
rect 5408 12180 5414 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 6362 12220 6368 12232
rect 6323 12192 6368 12220
rect 5445 12183 5503 12189
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 6779 12192 8309 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 6549 12155 6607 12161
rect 6549 12121 6561 12155
rect 6595 12152 6607 12155
rect 6595 12124 6776 12152
rect 6595 12121 6607 12124
rect 6549 12115 6607 12121
rect 6748 12096 6776 12124
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 3973 12087 4031 12093
rect 3973 12084 3985 12087
rect 3568 12056 3985 12084
rect 3568 12044 3574 12056
rect 3973 12053 3985 12056
rect 4019 12053 4031 12087
rect 5258 12084 5264 12096
rect 5219 12056 5264 12084
rect 3973 12047 4031 12053
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 6730 12044 6736 12096
rect 6788 12044 6794 12096
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 8570 12084 8576 12096
rect 8527 12056 8576 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 8570 12044 8576 12056
rect 8628 12044 8634 12096
rect 1104 11994 16995 12016
rect 1104 11942 4882 11994
rect 4934 11942 4946 11994
rect 4998 11942 5010 11994
rect 5062 11942 5074 11994
rect 5126 11942 5138 11994
rect 5190 11942 8815 11994
rect 8867 11942 8879 11994
rect 8931 11942 8943 11994
rect 8995 11942 9007 11994
rect 9059 11942 9071 11994
rect 9123 11942 12748 11994
rect 12800 11942 12812 11994
rect 12864 11942 12876 11994
rect 12928 11942 12940 11994
rect 12992 11942 13004 11994
rect 13056 11942 16681 11994
rect 16733 11942 16745 11994
rect 16797 11942 16809 11994
rect 16861 11942 16873 11994
rect 16925 11942 16937 11994
rect 16989 11942 16995 11994
rect 1104 11920 16995 11942
rect 3418 11880 3424 11892
rect 3379 11852 3424 11880
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 5077 11883 5135 11889
rect 5077 11880 5089 11883
rect 4304 11852 5089 11880
rect 4304 11840 4310 11852
rect 5077 11849 5089 11852
rect 5123 11849 5135 11883
rect 5258 11880 5264 11892
rect 5219 11852 5264 11880
rect 5077 11843 5135 11849
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 5350 11812 5356 11824
rect 3620 11784 5356 11812
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 3418 11744 3424 11756
rect 2363 11716 3424 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 3620 11753 3648 11784
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 6270 11812 6276 11824
rect 5592 11784 6276 11812
rect 5592 11772 5598 11784
rect 6270 11772 6276 11784
rect 6328 11812 6334 11824
rect 6328 11784 8892 11812
rect 6328 11772 6334 11784
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11713 3663 11747
rect 3878 11744 3884 11756
rect 3839 11716 3884 11744
rect 3605 11707 3663 11713
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 4062 11744 4068 11756
rect 4023 11716 4068 11744
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 5258 11747 5316 11753
rect 5258 11713 5270 11747
rect 5304 11744 5316 11747
rect 5442 11744 5448 11756
rect 5304 11716 5448 11744
rect 5304 11713 5316 11716
rect 5258 11707 5316 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 8570 11744 8576 11756
rect 8531 11716 8576 11744
rect 6549 11707 6607 11713
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 3896 11676 3924 11704
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 2648 11648 2693 11676
rect 3896 11648 5733 11676
rect 2648 11636 2654 11648
rect 5721 11645 5733 11648
rect 5767 11676 5779 11679
rect 5902 11676 5908 11688
rect 5767 11648 5908 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 6564 11608 6592 11707
rect 8570 11704 8576 11716
rect 8628 11704 8634 11756
rect 8864 11753 8892 11784
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 4764 11580 6592 11608
rect 4764 11568 4770 11580
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 4120 11512 5641 11540
rect 4120 11500 4126 11512
rect 5629 11509 5641 11512
rect 5675 11540 5687 11543
rect 5994 11540 6000 11552
rect 5675 11512 6000 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 5994 11500 6000 11512
rect 6052 11540 6058 11552
rect 6733 11543 6791 11549
rect 6733 11540 6745 11543
rect 6052 11512 6745 11540
rect 6052 11500 6058 11512
rect 6733 11509 6745 11512
rect 6779 11509 6791 11543
rect 9582 11540 9588 11552
rect 9543 11512 9588 11540
rect 6733 11503 6791 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 1104 11450 16836 11472
rect 1104 11398 2916 11450
rect 2968 11398 2980 11450
rect 3032 11398 3044 11450
rect 3096 11398 3108 11450
rect 3160 11398 3172 11450
rect 3224 11398 6849 11450
rect 6901 11398 6913 11450
rect 6965 11398 6977 11450
rect 7029 11398 7041 11450
rect 7093 11398 7105 11450
rect 7157 11398 10782 11450
rect 10834 11398 10846 11450
rect 10898 11398 10910 11450
rect 10962 11398 10974 11450
rect 11026 11398 11038 11450
rect 11090 11398 14715 11450
rect 14767 11398 14779 11450
rect 14831 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 16836 11450
rect 1104 11376 16836 11398
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 3326 11336 3332 11348
rect 2823 11308 3332 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 4055 11339 4113 11345
rect 4055 11336 4067 11339
rect 3476 11308 4067 11336
rect 3476 11296 3482 11308
rect 4055 11305 4067 11308
rect 4101 11336 4113 11339
rect 13354 11336 13360 11348
rect 4101 11308 13360 11336
rect 4101 11305 4113 11308
rect 4055 11299 4113 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 1854 11268 1860 11280
rect 1815 11240 1860 11268
rect 1854 11228 1860 11240
rect 1912 11228 1918 11280
rect 3237 11271 3295 11277
rect 3237 11237 3249 11271
rect 3283 11268 3295 11271
rect 3602 11268 3608 11280
rect 3283 11240 3608 11268
rect 3283 11237 3295 11240
rect 3237 11231 3295 11237
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 5537 11271 5595 11277
rect 5537 11237 5549 11271
rect 5583 11268 5595 11271
rect 5810 11268 5816 11280
rect 5583 11240 5816 11268
rect 5583 11237 5595 11240
rect 5537 11231 5595 11237
rect 5810 11228 5816 11240
rect 5868 11228 5874 11280
rect 5902 11228 5908 11280
rect 5960 11268 5966 11280
rect 5960 11240 6005 11268
rect 5960 11228 5966 11240
rect 5994 11200 6000 11212
rect 5955 11172 6000 11200
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 1670 11132 1676 11144
rect 1631 11104 1676 11132
rect 1670 11092 1676 11104
rect 1728 11092 1734 11144
rect 2406 11092 2412 11144
rect 2464 11132 2470 11144
rect 2593 11135 2651 11141
rect 2593 11132 2605 11135
rect 2464 11104 2605 11132
rect 2464 11092 2470 11104
rect 2593 11101 2605 11104
rect 2639 11101 2651 11135
rect 2593 11095 2651 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3510 11132 3516 11144
rect 3467 11104 3516 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4801 11135 4859 11141
rect 4801 11132 4813 11135
rect 4304 11104 4813 11132
rect 4304 11092 4310 11104
rect 4801 11101 4813 11104
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5626 11132 5632 11144
rect 5123 11104 5632 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 1688 11064 1716 11092
rect 2774 11064 2780 11076
rect 1688 11036 2780 11064
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 5736 11064 5764 11095
rect 7190 11064 7196 11076
rect 5736 11036 7196 11064
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 1104 10906 16995 10928
rect 1104 10854 4882 10906
rect 4934 10854 4946 10906
rect 4998 10854 5010 10906
rect 5062 10854 5074 10906
rect 5126 10854 5138 10906
rect 5190 10854 8815 10906
rect 8867 10854 8879 10906
rect 8931 10854 8943 10906
rect 8995 10854 9007 10906
rect 9059 10854 9071 10906
rect 9123 10854 12748 10906
rect 12800 10854 12812 10906
rect 12864 10854 12876 10906
rect 12928 10854 12940 10906
rect 12992 10854 13004 10906
rect 13056 10854 16681 10906
rect 16733 10854 16745 10906
rect 16797 10854 16809 10906
rect 16861 10854 16873 10906
rect 16925 10854 16937 10906
rect 16989 10854 16995 10906
rect 1104 10832 16995 10854
rect 2774 10792 2780 10804
rect 2735 10764 2780 10792
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 4157 10795 4215 10801
rect 4157 10761 4169 10795
rect 4203 10792 4215 10795
rect 4798 10792 4804 10804
rect 4203 10764 4804 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 5684 10764 6561 10792
rect 5684 10752 5690 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 6549 10755 6607 10761
rect 1854 10684 1860 10736
rect 1912 10724 1918 10736
rect 1949 10727 2007 10733
rect 1949 10724 1961 10727
rect 1912 10696 1961 10724
rect 1912 10684 1918 10696
rect 1949 10693 1961 10696
rect 1995 10693 2007 10727
rect 1949 10687 2007 10693
rect 5994 10684 6000 10736
rect 6052 10724 6058 10736
rect 6052 10696 6960 10724
rect 6052 10684 6058 10696
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10656 2191 10659
rect 2222 10656 2228 10668
rect 2179 10628 2228 10656
rect 2179 10625 2191 10628
rect 2133 10619 2191 10625
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 2363 10628 3709 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 3697 10625 3709 10628
rect 3743 10656 3755 10659
rect 3878 10656 3884 10668
rect 3743 10628 3884 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 4580 10628 5365 10656
rect 4580 10616 4586 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 6730 10656 6736 10668
rect 6691 10628 6736 10656
rect 5353 10619 5411 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 6932 10665 6960 10696
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 6840 10588 6868 10619
rect 9582 10588 9588 10600
rect 6840 10560 9588 10588
rect 3694 10480 3700 10532
rect 3752 10520 3758 10532
rect 6886 10520 6914 10560
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 3752 10492 6914 10520
rect 3752 10480 3758 10492
rect 3973 10455 4031 10461
rect 3973 10421 3985 10455
rect 4019 10452 4031 10455
rect 4062 10452 4068 10464
rect 4019 10424 4068 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 1104 10362 16836 10384
rect 1104 10310 2916 10362
rect 2968 10310 2980 10362
rect 3032 10310 3044 10362
rect 3096 10310 3108 10362
rect 3160 10310 3172 10362
rect 3224 10310 6849 10362
rect 6901 10310 6913 10362
rect 6965 10310 6977 10362
rect 7029 10310 7041 10362
rect 7093 10310 7105 10362
rect 7157 10310 10782 10362
rect 10834 10310 10846 10362
rect 10898 10310 10910 10362
rect 10962 10310 10974 10362
rect 11026 10310 11038 10362
rect 11090 10310 14715 10362
rect 14767 10310 14779 10362
rect 14831 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 16836 10362
rect 1104 10288 16836 10310
rect 1765 10251 1823 10257
rect 1765 10217 1777 10251
rect 1811 10248 1823 10251
rect 4154 10248 4160 10260
rect 1811 10220 4160 10248
rect 1811 10217 1823 10220
rect 1765 10211 1823 10217
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4304 10220 4353 10248
rect 4304 10208 4310 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 4522 10248 4528 10260
rect 4483 10220 4528 10248
rect 4341 10211 4399 10217
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 7101 10251 7159 10257
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7190 10248 7196 10260
rect 7147 10220 7196 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 2222 10140 2228 10192
rect 2280 10180 2286 10192
rect 3973 10183 4031 10189
rect 3973 10180 3985 10183
rect 2280 10152 3985 10180
rect 2280 10140 2286 10152
rect 3973 10149 3985 10152
rect 4019 10180 4031 10183
rect 6730 10180 6736 10192
rect 4019 10152 6736 10180
rect 4019 10149 4031 10152
rect 3973 10143 4031 10149
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 7374 10112 7380 10124
rect 7335 10084 7380 10112
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 1854 10044 1860 10056
rect 1815 10016 1860 10044
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 4341 9979 4399 9985
rect 4341 9945 4353 9979
rect 4387 9976 4399 9979
rect 4706 9976 4712 9988
rect 4387 9948 4712 9976
rect 4387 9945 4399 9948
rect 4341 9939 4399 9945
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 1104 9818 16995 9840
rect 1104 9766 4882 9818
rect 4934 9766 4946 9818
rect 4998 9766 5010 9818
rect 5062 9766 5074 9818
rect 5126 9766 5138 9818
rect 5190 9766 8815 9818
rect 8867 9766 8879 9818
rect 8931 9766 8943 9818
rect 8995 9766 9007 9818
rect 9059 9766 9071 9818
rect 9123 9766 12748 9818
rect 12800 9766 12812 9818
rect 12864 9766 12876 9818
rect 12928 9766 12940 9818
rect 12992 9766 13004 9818
rect 13056 9766 16681 9818
rect 16733 9766 16745 9818
rect 16797 9766 16809 9818
rect 16861 9766 16873 9818
rect 16925 9766 16937 9818
rect 16989 9766 16995 9818
rect 1104 9744 16995 9766
rect 2222 9568 2228 9580
rect 2183 9540 2228 9568
rect 2222 9528 2228 9540
rect 2280 9568 2286 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 2280 9540 4077 9568
rect 2280 9528 2286 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 4706 9500 4712 9512
rect 3835 9472 4712 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 2406 9432 2412 9444
rect 2367 9404 2412 9432
rect 2406 9392 2412 9404
rect 2464 9392 2470 9444
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 1912 9336 3525 9364
rect 1912 9324 1918 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3694 9364 3700 9376
rect 3655 9336 3700 9364
rect 3513 9327 3571 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 1104 9274 16836 9296
rect 1104 9222 2916 9274
rect 2968 9222 2980 9274
rect 3032 9222 3044 9274
rect 3096 9222 3108 9274
rect 3160 9222 3172 9274
rect 3224 9222 6849 9274
rect 6901 9222 6913 9274
rect 6965 9222 6977 9274
rect 7029 9222 7041 9274
rect 7093 9222 7105 9274
rect 7157 9222 10782 9274
rect 10834 9222 10846 9274
rect 10898 9222 10910 9274
rect 10962 9222 10974 9274
rect 11026 9222 11038 9274
rect 11090 9222 14715 9274
rect 14767 9222 14779 9274
rect 14831 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 16836 9274
rect 1104 9200 16836 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2590 9160 2596 9172
rect 2087 9132 2596 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 1104 8730 16995 8752
rect 1104 8678 4882 8730
rect 4934 8678 4946 8730
rect 4998 8678 5010 8730
rect 5062 8678 5074 8730
rect 5126 8678 5138 8730
rect 5190 8678 8815 8730
rect 8867 8678 8879 8730
rect 8931 8678 8943 8730
rect 8995 8678 9007 8730
rect 9059 8678 9071 8730
rect 9123 8678 12748 8730
rect 12800 8678 12812 8730
rect 12864 8678 12876 8730
rect 12928 8678 12940 8730
rect 12992 8678 13004 8730
rect 13056 8678 16681 8730
rect 16733 8678 16745 8730
rect 16797 8678 16809 8730
rect 16861 8678 16873 8730
rect 16925 8678 16937 8730
rect 16989 8678 16995 8730
rect 1104 8656 16995 8678
rect 1104 8186 16836 8208
rect 1104 8134 2916 8186
rect 2968 8134 2980 8186
rect 3032 8134 3044 8186
rect 3096 8134 3108 8186
rect 3160 8134 3172 8186
rect 3224 8134 6849 8186
rect 6901 8134 6913 8186
rect 6965 8134 6977 8186
rect 7029 8134 7041 8186
rect 7093 8134 7105 8186
rect 7157 8134 10782 8186
rect 10834 8134 10846 8186
rect 10898 8134 10910 8186
rect 10962 8134 10974 8186
rect 11026 8134 11038 8186
rect 11090 8134 14715 8186
rect 14767 8134 14779 8186
rect 14831 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 16836 8186
rect 1104 8112 16836 8134
rect 1104 7642 16995 7664
rect 1104 7590 4882 7642
rect 4934 7590 4946 7642
rect 4998 7590 5010 7642
rect 5062 7590 5074 7642
rect 5126 7590 5138 7642
rect 5190 7590 8815 7642
rect 8867 7590 8879 7642
rect 8931 7590 8943 7642
rect 8995 7590 9007 7642
rect 9059 7590 9071 7642
rect 9123 7590 12748 7642
rect 12800 7590 12812 7642
rect 12864 7590 12876 7642
rect 12928 7590 12940 7642
rect 12992 7590 13004 7642
rect 13056 7590 16681 7642
rect 16733 7590 16745 7642
rect 16797 7590 16809 7642
rect 16861 7590 16873 7642
rect 16925 7590 16937 7642
rect 16989 7590 16995 7642
rect 1104 7568 16995 7590
rect 1104 7098 16836 7120
rect 1104 7046 2916 7098
rect 2968 7046 2980 7098
rect 3032 7046 3044 7098
rect 3096 7046 3108 7098
rect 3160 7046 3172 7098
rect 3224 7046 6849 7098
rect 6901 7046 6913 7098
rect 6965 7046 6977 7098
rect 7029 7046 7041 7098
rect 7093 7046 7105 7098
rect 7157 7046 10782 7098
rect 10834 7046 10846 7098
rect 10898 7046 10910 7098
rect 10962 7046 10974 7098
rect 11026 7046 11038 7098
rect 11090 7046 14715 7098
rect 14767 7046 14779 7098
rect 14831 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 16836 7098
rect 1104 7024 16836 7046
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 1581 6783 1639 6789
rect 1581 6780 1593 6783
rect 1544 6752 1593 6780
rect 1544 6740 1550 6752
rect 1581 6749 1593 6752
rect 1627 6780 1639 6783
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 1627 6752 2237 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 2225 6749 2237 6752
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 4246 6712 4252 6724
rect 1780 6684 4252 6712
rect 1780 6653 1808 6684
rect 4246 6672 4252 6684
rect 4304 6672 4310 6724
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6613 1823 6647
rect 1765 6607 1823 6613
rect 1104 6554 16995 6576
rect 1104 6502 4882 6554
rect 4934 6502 4946 6554
rect 4998 6502 5010 6554
rect 5062 6502 5074 6554
rect 5126 6502 5138 6554
rect 5190 6502 8815 6554
rect 8867 6502 8879 6554
rect 8931 6502 8943 6554
rect 8995 6502 9007 6554
rect 9059 6502 9071 6554
rect 9123 6502 12748 6554
rect 12800 6502 12812 6554
rect 12864 6502 12876 6554
rect 12928 6502 12940 6554
rect 12992 6502 13004 6554
rect 13056 6502 16681 6554
rect 16733 6502 16745 6554
rect 16797 6502 16809 6554
rect 16861 6502 16873 6554
rect 16925 6502 16937 6554
rect 16989 6502 16995 6554
rect 1104 6480 16995 6502
rect 1104 6010 16836 6032
rect 1104 5958 2916 6010
rect 2968 5958 2980 6010
rect 3032 5958 3044 6010
rect 3096 5958 3108 6010
rect 3160 5958 3172 6010
rect 3224 5958 6849 6010
rect 6901 5958 6913 6010
rect 6965 5958 6977 6010
rect 7029 5958 7041 6010
rect 7093 5958 7105 6010
rect 7157 5958 10782 6010
rect 10834 5958 10846 6010
rect 10898 5958 10910 6010
rect 10962 5958 10974 6010
rect 11026 5958 11038 6010
rect 11090 5958 14715 6010
rect 14767 5958 14779 6010
rect 14831 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 16836 6010
rect 1104 5936 16836 5958
rect 1104 5466 16995 5488
rect 1104 5414 4882 5466
rect 4934 5414 4946 5466
rect 4998 5414 5010 5466
rect 5062 5414 5074 5466
rect 5126 5414 5138 5466
rect 5190 5414 8815 5466
rect 8867 5414 8879 5466
rect 8931 5414 8943 5466
rect 8995 5414 9007 5466
rect 9059 5414 9071 5466
rect 9123 5414 12748 5466
rect 12800 5414 12812 5466
rect 12864 5414 12876 5466
rect 12928 5414 12940 5466
rect 12992 5414 13004 5466
rect 13056 5414 16681 5466
rect 16733 5414 16745 5466
rect 16797 5414 16809 5466
rect 16861 5414 16873 5466
rect 16925 5414 16937 5466
rect 16989 5414 16995 5466
rect 1104 5392 16995 5414
rect 1104 4922 16836 4944
rect 1104 4870 2916 4922
rect 2968 4870 2980 4922
rect 3032 4870 3044 4922
rect 3096 4870 3108 4922
rect 3160 4870 3172 4922
rect 3224 4870 6849 4922
rect 6901 4870 6913 4922
rect 6965 4870 6977 4922
rect 7029 4870 7041 4922
rect 7093 4870 7105 4922
rect 7157 4870 10782 4922
rect 10834 4870 10846 4922
rect 10898 4870 10910 4922
rect 10962 4870 10974 4922
rect 11026 4870 11038 4922
rect 11090 4870 14715 4922
rect 14767 4870 14779 4922
rect 14831 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 16836 4922
rect 1104 4848 16836 4870
rect 1104 4378 16995 4400
rect 1104 4326 4882 4378
rect 4934 4326 4946 4378
rect 4998 4326 5010 4378
rect 5062 4326 5074 4378
rect 5126 4326 5138 4378
rect 5190 4326 8815 4378
rect 8867 4326 8879 4378
rect 8931 4326 8943 4378
rect 8995 4326 9007 4378
rect 9059 4326 9071 4378
rect 9123 4326 12748 4378
rect 12800 4326 12812 4378
rect 12864 4326 12876 4378
rect 12928 4326 12940 4378
rect 12992 4326 13004 4378
rect 13056 4326 16681 4378
rect 16733 4326 16745 4378
rect 16797 4326 16809 4378
rect 16861 4326 16873 4378
rect 16925 4326 16937 4378
rect 16989 4326 16995 4378
rect 1104 4304 16995 4326
rect 1104 3834 16836 3856
rect 1104 3782 2916 3834
rect 2968 3782 2980 3834
rect 3032 3782 3044 3834
rect 3096 3782 3108 3834
rect 3160 3782 3172 3834
rect 3224 3782 6849 3834
rect 6901 3782 6913 3834
rect 6965 3782 6977 3834
rect 7029 3782 7041 3834
rect 7093 3782 7105 3834
rect 7157 3782 10782 3834
rect 10834 3782 10846 3834
rect 10898 3782 10910 3834
rect 10962 3782 10974 3834
rect 11026 3782 11038 3834
rect 11090 3782 14715 3834
rect 14767 3782 14779 3834
rect 14831 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 16836 3834
rect 1104 3760 16836 3782
rect 1104 3290 16995 3312
rect 1104 3238 4882 3290
rect 4934 3238 4946 3290
rect 4998 3238 5010 3290
rect 5062 3238 5074 3290
rect 5126 3238 5138 3290
rect 5190 3238 8815 3290
rect 8867 3238 8879 3290
rect 8931 3238 8943 3290
rect 8995 3238 9007 3290
rect 9059 3238 9071 3290
rect 9123 3238 12748 3290
rect 12800 3238 12812 3290
rect 12864 3238 12876 3290
rect 12928 3238 12940 3290
rect 12992 3238 13004 3290
rect 13056 3238 16681 3290
rect 16733 3238 16745 3290
rect 16797 3238 16809 3290
rect 16861 3238 16873 3290
rect 16925 3238 16937 3290
rect 16989 3238 16995 3290
rect 1104 3216 16995 3238
rect 1104 2746 16836 2768
rect 1104 2694 2916 2746
rect 2968 2694 2980 2746
rect 3032 2694 3044 2746
rect 3096 2694 3108 2746
rect 3160 2694 3172 2746
rect 3224 2694 6849 2746
rect 6901 2694 6913 2746
rect 6965 2694 6977 2746
rect 7029 2694 7041 2746
rect 7093 2694 7105 2746
rect 7157 2694 10782 2746
rect 10834 2694 10846 2746
rect 10898 2694 10910 2746
rect 10962 2694 10974 2746
rect 11026 2694 11038 2746
rect 11090 2694 14715 2746
rect 14767 2694 14779 2746
rect 14831 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 16836 2746
rect 1104 2672 16836 2694
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 1104 2202 16995 2224
rect 1104 2150 4882 2202
rect 4934 2150 4946 2202
rect 4998 2150 5010 2202
rect 5062 2150 5074 2202
rect 5126 2150 5138 2202
rect 5190 2150 8815 2202
rect 8867 2150 8879 2202
rect 8931 2150 8943 2202
rect 8995 2150 9007 2202
rect 9059 2150 9071 2202
rect 9123 2150 12748 2202
rect 12800 2150 12812 2202
rect 12864 2150 12876 2202
rect 12928 2150 12940 2202
rect 12992 2150 13004 2202
rect 13056 2150 16681 2202
rect 16733 2150 16745 2202
rect 16797 2150 16809 2202
rect 16861 2150 16873 2202
rect 16925 2150 16937 2202
rect 16989 2150 16995 2202
rect 1104 2128 16995 2150
<< via1 >>
rect 2916 15750 2968 15802
rect 2980 15750 3032 15802
rect 3044 15750 3096 15802
rect 3108 15750 3160 15802
rect 3172 15750 3224 15802
rect 6849 15750 6901 15802
rect 6913 15750 6965 15802
rect 6977 15750 7029 15802
rect 7041 15750 7093 15802
rect 7105 15750 7157 15802
rect 10782 15750 10834 15802
rect 10846 15750 10898 15802
rect 10910 15750 10962 15802
rect 10974 15750 11026 15802
rect 11038 15750 11090 15802
rect 14715 15750 14767 15802
rect 14779 15750 14831 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 1584 15648 1636 15700
rect 4528 15648 4580 15700
rect 7472 15648 7524 15700
rect 10692 15691 10744 15700
rect 10692 15657 10701 15691
rect 10701 15657 10735 15691
rect 10735 15657 10744 15691
rect 10692 15648 10744 15657
rect 16212 15691 16264 15700
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 3792 15580 3844 15632
rect 2044 15512 2096 15564
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 3700 15376 3752 15428
rect 3240 15308 3292 15360
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 6000 15487 6052 15496
rect 6000 15453 6009 15487
rect 6009 15453 6043 15487
rect 6043 15453 6052 15487
rect 6000 15444 6052 15453
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 8300 15444 8352 15496
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 4882 15206 4934 15258
rect 4946 15206 4998 15258
rect 5010 15206 5062 15258
rect 5074 15206 5126 15258
rect 5138 15206 5190 15258
rect 8815 15206 8867 15258
rect 8879 15206 8931 15258
rect 8943 15206 8995 15258
rect 9007 15206 9059 15258
rect 9071 15206 9123 15258
rect 12748 15206 12800 15258
rect 12812 15206 12864 15258
rect 12876 15206 12928 15258
rect 12940 15206 12992 15258
rect 13004 15206 13056 15258
rect 16681 15206 16733 15258
rect 16745 15206 16797 15258
rect 16809 15206 16861 15258
rect 16873 15206 16925 15258
rect 16937 15206 16989 15258
rect 2044 15104 2096 15156
rect 6552 15104 6604 15156
rect 8300 15104 8352 15156
rect 3608 15036 3660 15088
rect 6276 15036 6328 15088
rect 5448 14968 5500 15020
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 6552 14968 6604 15020
rect 2688 14900 2740 14952
rect 3332 14943 3384 14952
rect 3332 14909 3341 14943
rect 3341 14909 3375 14943
rect 3375 14909 3384 14943
rect 3332 14900 3384 14909
rect 2780 14764 2832 14816
rect 2916 14662 2968 14714
rect 2980 14662 3032 14714
rect 3044 14662 3096 14714
rect 3108 14662 3160 14714
rect 3172 14662 3224 14714
rect 6849 14662 6901 14714
rect 6913 14662 6965 14714
rect 6977 14662 7029 14714
rect 7041 14662 7093 14714
rect 7105 14662 7157 14714
rect 10782 14662 10834 14714
rect 10846 14662 10898 14714
rect 10910 14662 10962 14714
rect 10974 14662 11026 14714
rect 11038 14662 11090 14714
rect 14715 14662 14767 14714
rect 14779 14662 14831 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 5816 14560 5868 14612
rect 6828 14560 6880 14612
rect 7564 14560 7616 14612
rect 5816 14424 5868 14476
rect 2780 14356 2832 14408
rect 3884 14356 3936 14408
rect 6552 14399 6604 14408
rect 6552 14365 6561 14399
rect 6561 14365 6595 14399
rect 6595 14365 6604 14399
rect 6552 14356 6604 14365
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 2136 14263 2188 14272
rect 2136 14229 2145 14263
rect 2145 14229 2179 14263
rect 2179 14229 2188 14263
rect 2136 14220 2188 14229
rect 3700 14220 3752 14272
rect 6644 14220 6696 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 4882 14118 4934 14170
rect 4946 14118 4998 14170
rect 5010 14118 5062 14170
rect 5074 14118 5126 14170
rect 5138 14118 5190 14170
rect 8815 14118 8867 14170
rect 8879 14118 8931 14170
rect 8943 14118 8995 14170
rect 9007 14118 9059 14170
rect 9071 14118 9123 14170
rect 12748 14118 12800 14170
rect 12812 14118 12864 14170
rect 12876 14118 12928 14170
rect 12940 14118 12992 14170
rect 13004 14118 13056 14170
rect 16681 14118 16733 14170
rect 16745 14118 16797 14170
rect 16809 14118 16861 14170
rect 16873 14118 16925 14170
rect 16937 14118 16989 14170
rect 1584 14016 1636 14068
rect 2688 14016 2740 14068
rect 6736 14016 6788 14068
rect 4160 13948 4212 14000
rect 5724 13948 5776 14000
rect 6000 13991 6052 14000
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 5632 13923 5684 13932
rect 5632 13889 5641 13923
rect 5641 13889 5675 13923
rect 5675 13889 5684 13923
rect 6000 13957 6009 13991
rect 6009 13957 6043 13991
rect 6043 13957 6052 13991
rect 6000 13948 6052 13957
rect 6644 13948 6696 14000
rect 5632 13880 5684 13889
rect 3424 13855 3476 13864
rect 2228 13676 2280 13728
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 3884 13676 3936 13728
rect 5264 13676 5316 13728
rect 5448 13676 5500 13728
rect 7196 13923 7248 13932
rect 7196 13889 7205 13923
rect 7205 13889 7239 13923
rect 7239 13889 7248 13923
rect 7196 13880 7248 13889
rect 7288 13812 7340 13864
rect 2916 13574 2968 13626
rect 2980 13574 3032 13626
rect 3044 13574 3096 13626
rect 3108 13574 3160 13626
rect 3172 13574 3224 13626
rect 6849 13574 6901 13626
rect 6913 13574 6965 13626
rect 6977 13574 7029 13626
rect 7041 13574 7093 13626
rect 7105 13574 7157 13626
rect 10782 13574 10834 13626
rect 10846 13574 10898 13626
rect 10910 13574 10962 13626
rect 10974 13574 11026 13626
rect 11038 13574 11090 13626
rect 14715 13574 14767 13626
rect 14779 13574 14831 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 4436 13472 4488 13524
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 7748 13472 7800 13524
rect 4620 13336 4672 13388
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 7196 13379 7248 13388
rect 5724 13336 5776 13345
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 3884 13268 3936 13320
rect 6184 13311 6236 13320
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 6184 13268 6236 13277
rect 6276 13268 6328 13320
rect 6552 13268 6604 13320
rect 6644 13268 6696 13320
rect 3240 13200 3292 13252
rect 4252 13243 4304 13252
rect 4252 13209 4261 13243
rect 4261 13209 4295 13243
rect 4295 13209 4304 13243
rect 4252 13200 4304 13209
rect 3700 13132 3752 13184
rect 4882 13030 4934 13082
rect 4946 13030 4998 13082
rect 5010 13030 5062 13082
rect 5074 13030 5126 13082
rect 5138 13030 5190 13082
rect 8815 13030 8867 13082
rect 8879 13030 8931 13082
rect 8943 13030 8995 13082
rect 9007 13030 9059 13082
rect 9071 13030 9123 13082
rect 12748 13030 12800 13082
rect 12812 13030 12864 13082
rect 12876 13030 12928 13082
rect 12940 13030 12992 13082
rect 13004 13030 13056 13082
rect 16681 13030 16733 13082
rect 16745 13030 16797 13082
rect 16809 13030 16861 13082
rect 16873 13030 16925 13082
rect 16937 13030 16989 13082
rect 3700 12928 3752 12980
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 5540 12928 5592 12980
rect 2136 12860 2188 12912
rect 2596 12903 2648 12912
rect 2596 12869 2605 12903
rect 2605 12869 2639 12903
rect 2639 12869 2648 12903
rect 2596 12860 2648 12869
rect 1860 12792 1912 12844
rect 2412 12792 2464 12844
rect 6184 12860 6236 12912
rect 4620 12792 4672 12844
rect 4804 12792 4856 12844
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5632 12792 5684 12844
rect 6644 12792 6696 12844
rect 5724 12724 5776 12776
rect 7288 12792 7340 12844
rect 7472 12724 7524 12776
rect 6368 12588 6420 12640
rect 7196 12588 7248 12640
rect 2916 12486 2968 12538
rect 2980 12486 3032 12538
rect 3044 12486 3096 12538
rect 3108 12486 3160 12538
rect 3172 12486 3224 12538
rect 6849 12486 6901 12538
rect 6913 12486 6965 12538
rect 6977 12486 7029 12538
rect 7041 12486 7093 12538
rect 7105 12486 7157 12538
rect 10782 12486 10834 12538
rect 10846 12486 10898 12538
rect 10910 12486 10962 12538
rect 10974 12486 11026 12538
rect 11038 12486 11090 12538
rect 14715 12486 14767 12538
rect 14779 12486 14831 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 4620 12427 4672 12436
rect 4620 12393 4629 12427
rect 4629 12393 4663 12427
rect 4663 12393 4672 12427
rect 4620 12384 4672 12393
rect 1584 12291 1636 12300
rect 1584 12257 1593 12291
rect 1593 12257 1627 12291
rect 1627 12257 1636 12291
rect 1584 12248 1636 12257
rect 5632 12248 5684 12300
rect 5724 12248 5776 12300
rect 2596 12180 2648 12232
rect 4068 12180 4120 12232
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 5356 12180 5408 12232
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 3516 12044 3568 12096
rect 5264 12087 5316 12096
rect 5264 12053 5273 12087
rect 5273 12053 5307 12087
rect 5307 12053 5316 12087
rect 5264 12044 5316 12053
rect 6736 12044 6788 12096
rect 8576 12044 8628 12096
rect 4882 11942 4934 11994
rect 4946 11942 4998 11994
rect 5010 11942 5062 11994
rect 5074 11942 5126 11994
rect 5138 11942 5190 11994
rect 8815 11942 8867 11994
rect 8879 11942 8931 11994
rect 8943 11942 8995 11994
rect 9007 11942 9059 11994
rect 9071 11942 9123 11994
rect 12748 11942 12800 11994
rect 12812 11942 12864 11994
rect 12876 11942 12928 11994
rect 12940 11942 12992 11994
rect 13004 11942 13056 11994
rect 16681 11942 16733 11994
rect 16745 11942 16797 11994
rect 16809 11942 16861 11994
rect 16873 11942 16925 11994
rect 16937 11942 16989 11994
rect 3424 11883 3476 11892
rect 3424 11849 3433 11883
rect 3433 11849 3467 11883
rect 3467 11849 3476 11883
rect 3424 11840 3476 11849
rect 4252 11840 4304 11892
rect 5264 11883 5316 11892
rect 5264 11849 5273 11883
rect 5273 11849 5307 11883
rect 5307 11849 5316 11883
rect 5264 11840 5316 11849
rect 3424 11704 3476 11756
rect 5356 11772 5408 11824
rect 5540 11772 5592 11824
rect 6276 11772 6328 11824
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 5448 11704 5500 11756
rect 8576 11747 8628 11756
rect 2596 11679 2648 11688
rect 2596 11645 2605 11679
rect 2605 11645 2639 11679
rect 2639 11645 2648 11679
rect 2596 11636 2648 11645
rect 5908 11636 5960 11688
rect 4712 11568 4764 11620
rect 8576 11713 8585 11747
rect 8585 11713 8619 11747
rect 8619 11713 8628 11747
rect 8576 11704 8628 11713
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 4068 11500 4120 11552
rect 6000 11500 6052 11552
rect 9588 11543 9640 11552
rect 9588 11509 9597 11543
rect 9597 11509 9631 11543
rect 9631 11509 9640 11543
rect 9588 11500 9640 11509
rect 2916 11398 2968 11450
rect 2980 11398 3032 11450
rect 3044 11398 3096 11450
rect 3108 11398 3160 11450
rect 3172 11398 3224 11450
rect 6849 11398 6901 11450
rect 6913 11398 6965 11450
rect 6977 11398 7029 11450
rect 7041 11398 7093 11450
rect 7105 11398 7157 11450
rect 10782 11398 10834 11450
rect 10846 11398 10898 11450
rect 10910 11398 10962 11450
rect 10974 11398 11026 11450
rect 11038 11398 11090 11450
rect 14715 11398 14767 11450
rect 14779 11398 14831 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 3332 11296 3384 11348
rect 3424 11296 3476 11348
rect 13360 11296 13412 11348
rect 1860 11271 1912 11280
rect 1860 11237 1869 11271
rect 1869 11237 1903 11271
rect 1903 11237 1912 11271
rect 1860 11228 1912 11237
rect 3608 11228 3660 11280
rect 5816 11228 5868 11280
rect 5908 11271 5960 11280
rect 5908 11237 5917 11271
rect 5917 11237 5951 11271
rect 5951 11237 5960 11271
rect 5908 11228 5960 11237
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 2412 11092 2464 11144
rect 3516 11092 3568 11144
rect 4252 11092 4304 11144
rect 5632 11092 5684 11144
rect 2780 11024 2832 11076
rect 7196 11024 7248 11076
rect 4882 10854 4934 10906
rect 4946 10854 4998 10906
rect 5010 10854 5062 10906
rect 5074 10854 5126 10906
rect 5138 10854 5190 10906
rect 8815 10854 8867 10906
rect 8879 10854 8931 10906
rect 8943 10854 8995 10906
rect 9007 10854 9059 10906
rect 9071 10854 9123 10906
rect 12748 10854 12800 10906
rect 12812 10854 12864 10906
rect 12876 10854 12928 10906
rect 12940 10854 12992 10906
rect 13004 10854 13056 10906
rect 16681 10854 16733 10906
rect 16745 10854 16797 10906
rect 16809 10854 16861 10906
rect 16873 10854 16925 10906
rect 16937 10854 16989 10906
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 2780 10752 2832 10761
rect 4804 10752 4856 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 5632 10752 5684 10804
rect 1860 10684 1912 10736
rect 6000 10684 6052 10736
rect 2228 10616 2280 10668
rect 3884 10616 3936 10668
rect 4528 10616 4580 10668
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 3700 10480 3752 10532
rect 9588 10548 9640 10600
rect 4068 10412 4120 10464
rect 2916 10310 2968 10362
rect 2980 10310 3032 10362
rect 3044 10310 3096 10362
rect 3108 10310 3160 10362
rect 3172 10310 3224 10362
rect 6849 10310 6901 10362
rect 6913 10310 6965 10362
rect 6977 10310 7029 10362
rect 7041 10310 7093 10362
rect 7105 10310 7157 10362
rect 10782 10310 10834 10362
rect 10846 10310 10898 10362
rect 10910 10310 10962 10362
rect 10974 10310 11026 10362
rect 11038 10310 11090 10362
rect 14715 10310 14767 10362
rect 14779 10310 14831 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 4160 10208 4212 10260
rect 4252 10208 4304 10260
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 7196 10208 7248 10260
rect 2228 10140 2280 10192
rect 6736 10140 6788 10192
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 4712 9936 4764 9988
rect 4882 9766 4934 9818
rect 4946 9766 4998 9818
rect 5010 9766 5062 9818
rect 5074 9766 5126 9818
rect 5138 9766 5190 9818
rect 8815 9766 8867 9818
rect 8879 9766 8931 9818
rect 8943 9766 8995 9818
rect 9007 9766 9059 9818
rect 9071 9766 9123 9818
rect 12748 9766 12800 9818
rect 12812 9766 12864 9818
rect 12876 9766 12928 9818
rect 12940 9766 12992 9818
rect 13004 9766 13056 9818
rect 16681 9766 16733 9818
rect 16745 9766 16797 9818
rect 16809 9766 16861 9818
rect 16873 9766 16925 9818
rect 16937 9766 16989 9818
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 4712 9460 4764 9512
rect 2412 9435 2464 9444
rect 2412 9401 2421 9435
rect 2421 9401 2455 9435
rect 2455 9401 2464 9435
rect 2412 9392 2464 9401
rect 1860 9324 1912 9376
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 2916 9222 2968 9274
rect 2980 9222 3032 9274
rect 3044 9222 3096 9274
rect 3108 9222 3160 9274
rect 3172 9222 3224 9274
rect 6849 9222 6901 9274
rect 6913 9222 6965 9274
rect 6977 9222 7029 9274
rect 7041 9222 7093 9274
rect 7105 9222 7157 9274
rect 10782 9222 10834 9274
rect 10846 9222 10898 9274
rect 10910 9222 10962 9274
rect 10974 9222 11026 9274
rect 11038 9222 11090 9274
rect 14715 9222 14767 9274
rect 14779 9222 14831 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 2596 9120 2648 9172
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 4882 8678 4934 8730
rect 4946 8678 4998 8730
rect 5010 8678 5062 8730
rect 5074 8678 5126 8730
rect 5138 8678 5190 8730
rect 8815 8678 8867 8730
rect 8879 8678 8931 8730
rect 8943 8678 8995 8730
rect 9007 8678 9059 8730
rect 9071 8678 9123 8730
rect 12748 8678 12800 8730
rect 12812 8678 12864 8730
rect 12876 8678 12928 8730
rect 12940 8678 12992 8730
rect 13004 8678 13056 8730
rect 16681 8678 16733 8730
rect 16745 8678 16797 8730
rect 16809 8678 16861 8730
rect 16873 8678 16925 8730
rect 16937 8678 16989 8730
rect 2916 8134 2968 8186
rect 2980 8134 3032 8186
rect 3044 8134 3096 8186
rect 3108 8134 3160 8186
rect 3172 8134 3224 8186
rect 6849 8134 6901 8186
rect 6913 8134 6965 8186
rect 6977 8134 7029 8186
rect 7041 8134 7093 8186
rect 7105 8134 7157 8186
rect 10782 8134 10834 8186
rect 10846 8134 10898 8186
rect 10910 8134 10962 8186
rect 10974 8134 11026 8186
rect 11038 8134 11090 8186
rect 14715 8134 14767 8186
rect 14779 8134 14831 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 4882 7590 4934 7642
rect 4946 7590 4998 7642
rect 5010 7590 5062 7642
rect 5074 7590 5126 7642
rect 5138 7590 5190 7642
rect 8815 7590 8867 7642
rect 8879 7590 8931 7642
rect 8943 7590 8995 7642
rect 9007 7590 9059 7642
rect 9071 7590 9123 7642
rect 12748 7590 12800 7642
rect 12812 7590 12864 7642
rect 12876 7590 12928 7642
rect 12940 7590 12992 7642
rect 13004 7590 13056 7642
rect 16681 7590 16733 7642
rect 16745 7590 16797 7642
rect 16809 7590 16861 7642
rect 16873 7590 16925 7642
rect 16937 7590 16989 7642
rect 2916 7046 2968 7098
rect 2980 7046 3032 7098
rect 3044 7046 3096 7098
rect 3108 7046 3160 7098
rect 3172 7046 3224 7098
rect 6849 7046 6901 7098
rect 6913 7046 6965 7098
rect 6977 7046 7029 7098
rect 7041 7046 7093 7098
rect 7105 7046 7157 7098
rect 10782 7046 10834 7098
rect 10846 7046 10898 7098
rect 10910 7046 10962 7098
rect 10974 7046 11026 7098
rect 11038 7046 11090 7098
rect 14715 7046 14767 7098
rect 14779 7046 14831 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 1492 6740 1544 6792
rect 4252 6672 4304 6724
rect 4882 6502 4934 6554
rect 4946 6502 4998 6554
rect 5010 6502 5062 6554
rect 5074 6502 5126 6554
rect 5138 6502 5190 6554
rect 8815 6502 8867 6554
rect 8879 6502 8931 6554
rect 8943 6502 8995 6554
rect 9007 6502 9059 6554
rect 9071 6502 9123 6554
rect 12748 6502 12800 6554
rect 12812 6502 12864 6554
rect 12876 6502 12928 6554
rect 12940 6502 12992 6554
rect 13004 6502 13056 6554
rect 16681 6502 16733 6554
rect 16745 6502 16797 6554
rect 16809 6502 16861 6554
rect 16873 6502 16925 6554
rect 16937 6502 16989 6554
rect 2916 5958 2968 6010
rect 2980 5958 3032 6010
rect 3044 5958 3096 6010
rect 3108 5958 3160 6010
rect 3172 5958 3224 6010
rect 6849 5958 6901 6010
rect 6913 5958 6965 6010
rect 6977 5958 7029 6010
rect 7041 5958 7093 6010
rect 7105 5958 7157 6010
rect 10782 5958 10834 6010
rect 10846 5958 10898 6010
rect 10910 5958 10962 6010
rect 10974 5958 11026 6010
rect 11038 5958 11090 6010
rect 14715 5958 14767 6010
rect 14779 5958 14831 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 4882 5414 4934 5466
rect 4946 5414 4998 5466
rect 5010 5414 5062 5466
rect 5074 5414 5126 5466
rect 5138 5414 5190 5466
rect 8815 5414 8867 5466
rect 8879 5414 8931 5466
rect 8943 5414 8995 5466
rect 9007 5414 9059 5466
rect 9071 5414 9123 5466
rect 12748 5414 12800 5466
rect 12812 5414 12864 5466
rect 12876 5414 12928 5466
rect 12940 5414 12992 5466
rect 13004 5414 13056 5466
rect 16681 5414 16733 5466
rect 16745 5414 16797 5466
rect 16809 5414 16861 5466
rect 16873 5414 16925 5466
rect 16937 5414 16989 5466
rect 2916 4870 2968 4922
rect 2980 4870 3032 4922
rect 3044 4870 3096 4922
rect 3108 4870 3160 4922
rect 3172 4870 3224 4922
rect 6849 4870 6901 4922
rect 6913 4870 6965 4922
rect 6977 4870 7029 4922
rect 7041 4870 7093 4922
rect 7105 4870 7157 4922
rect 10782 4870 10834 4922
rect 10846 4870 10898 4922
rect 10910 4870 10962 4922
rect 10974 4870 11026 4922
rect 11038 4870 11090 4922
rect 14715 4870 14767 4922
rect 14779 4870 14831 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 4882 4326 4934 4378
rect 4946 4326 4998 4378
rect 5010 4326 5062 4378
rect 5074 4326 5126 4378
rect 5138 4326 5190 4378
rect 8815 4326 8867 4378
rect 8879 4326 8931 4378
rect 8943 4326 8995 4378
rect 9007 4326 9059 4378
rect 9071 4326 9123 4378
rect 12748 4326 12800 4378
rect 12812 4326 12864 4378
rect 12876 4326 12928 4378
rect 12940 4326 12992 4378
rect 13004 4326 13056 4378
rect 16681 4326 16733 4378
rect 16745 4326 16797 4378
rect 16809 4326 16861 4378
rect 16873 4326 16925 4378
rect 16937 4326 16989 4378
rect 2916 3782 2968 3834
rect 2980 3782 3032 3834
rect 3044 3782 3096 3834
rect 3108 3782 3160 3834
rect 3172 3782 3224 3834
rect 6849 3782 6901 3834
rect 6913 3782 6965 3834
rect 6977 3782 7029 3834
rect 7041 3782 7093 3834
rect 7105 3782 7157 3834
rect 10782 3782 10834 3834
rect 10846 3782 10898 3834
rect 10910 3782 10962 3834
rect 10974 3782 11026 3834
rect 11038 3782 11090 3834
rect 14715 3782 14767 3834
rect 14779 3782 14831 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 4882 3238 4934 3290
rect 4946 3238 4998 3290
rect 5010 3238 5062 3290
rect 5074 3238 5126 3290
rect 5138 3238 5190 3290
rect 8815 3238 8867 3290
rect 8879 3238 8931 3290
rect 8943 3238 8995 3290
rect 9007 3238 9059 3290
rect 9071 3238 9123 3290
rect 12748 3238 12800 3290
rect 12812 3238 12864 3290
rect 12876 3238 12928 3290
rect 12940 3238 12992 3290
rect 13004 3238 13056 3290
rect 16681 3238 16733 3290
rect 16745 3238 16797 3290
rect 16809 3238 16861 3290
rect 16873 3238 16925 3290
rect 16937 3238 16989 3290
rect 2916 2694 2968 2746
rect 2980 2694 3032 2746
rect 3044 2694 3096 2746
rect 3108 2694 3160 2746
rect 3172 2694 3224 2746
rect 6849 2694 6901 2746
rect 6913 2694 6965 2746
rect 6977 2694 7029 2746
rect 7041 2694 7093 2746
rect 7105 2694 7157 2746
rect 10782 2694 10834 2746
rect 10846 2694 10898 2746
rect 10910 2694 10962 2746
rect 10974 2694 11026 2746
rect 11038 2694 11090 2746
rect 14715 2694 14767 2746
rect 14779 2694 14831 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 4882 2150 4934 2202
rect 4946 2150 4998 2202
rect 5010 2150 5062 2202
rect 5074 2150 5126 2202
rect 5138 2150 5190 2202
rect 8815 2150 8867 2202
rect 8879 2150 8931 2202
rect 8943 2150 8995 2202
rect 9007 2150 9059 2202
rect 9071 2150 9123 2202
rect 12748 2150 12800 2202
rect 12812 2150 12864 2202
rect 12876 2150 12928 2202
rect 12940 2150 12992 2202
rect 13004 2150 13056 2202
rect 16681 2150 16733 2202
rect 16745 2150 16797 2202
rect 16809 2150 16861 2202
rect 16873 2150 16925 2202
rect 16937 2150 16989 2202
<< metal2 >>
rect 1582 17200 1638 18000
rect 4526 17200 4582 18000
rect 7470 17200 7526 18000
rect 10414 17354 10470 18000
rect 10414 17326 10732 17354
rect 10414 17200 10470 17326
rect 1596 15706 1624 17200
rect 2916 15804 3224 15813
rect 2916 15802 2922 15804
rect 2978 15802 3002 15804
rect 3058 15802 3082 15804
rect 3138 15802 3162 15804
rect 3218 15802 3224 15804
rect 2978 15750 2980 15802
rect 3160 15750 3162 15802
rect 2916 15748 2922 15750
rect 2978 15748 3002 15750
rect 3058 15748 3082 15750
rect 3138 15748 3162 15750
rect 3218 15748 3224 15750
rect 2778 15736 2834 15745
rect 2916 15739 3224 15748
rect 1584 15700 1636 15706
rect 4540 15706 4568 17200
rect 6849 15804 7157 15813
rect 6849 15802 6855 15804
rect 6911 15802 6935 15804
rect 6991 15802 7015 15804
rect 7071 15802 7095 15804
rect 7151 15802 7157 15804
rect 6911 15750 6913 15802
rect 7093 15750 7095 15802
rect 6849 15748 6855 15750
rect 6911 15748 6935 15750
rect 6991 15748 7015 15750
rect 7071 15748 7095 15750
rect 7151 15748 7157 15750
rect 6849 15739 7157 15748
rect 7484 15706 7512 17200
rect 10704 15706 10732 17326
rect 13358 17200 13414 18000
rect 16302 17354 16358 18000
rect 16224 17326 16358 17354
rect 10782 15804 11090 15813
rect 10782 15802 10788 15804
rect 10844 15802 10868 15804
rect 10924 15802 10948 15804
rect 11004 15802 11028 15804
rect 11084 15802 11090 15804
rect 10844 15750 10846 15802
rect 11026 15750 11028 15802
rect 10782 15748 10788 15750
rect 10844 15748 10868 15750
rect 10924 15748 10948 15750
rect 11004 15748 11028 15750
rect 11084 15748 11090 15750
rect 10782 15739 11090 15748
rect 2778 15671 2834 15680
rect 4528 15700 4580 15706
rect 1584 15642 1636 15648
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2056 15162 2084 15506
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1596 13394 1624 14010
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 12306 1624 13330
rect 2148 12918 2176 14214
rect 2226 13968 2282 13977
rect 2226 13903 2228 13912
rect 2280 13903 2282 13912
rect 2228 13874 2280 13880
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1492 6792 1544 6798
rect 1490 6760 1492 6769
rect 1544 6760 1546 6769
rect 1490 6695 1546 6704
rect 1596 2446 1624 11494
rect 1872 11286 1900 12786
rect 1860 11280 1912 11286
rect 1674 11248 1730 11257
rect 1860 11222 1912 11228
rect 1674 11183 1730 11192
rect 1688 11150 1716 11183
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1872 10742 1900 11222
rect 1860 10736 1912 10742
rect 1860 10678 1912 10684
rect 1872 10062 1900 10678
rect 2240 10674 2268 13670
rect 2424 12850 2452 15438
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2700 14074 2728 14894
rect 2792 14822 2820 15671
rect 4528 15642 4580 15648
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3700 15428 3752 15434
rect 3700 15370 3752 15376
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 14414 2820 14758
rect 2916 14716 3224 14725
rect 2916 14714 2922 14716
rect 2978 14714 3002 14716
rect 3058 14714 3082 14716
rect 3138 14714 3162 14716
rect 3218 14714 3224 14716
rect 2978 14662 2980 14714
rect 3160 14662 3162 14714
rect 2916 14660 2922 14662
rect 2978 14660 3002 14662
rect 3058 14660 3082 14662
rect 3138 14660 3162 14662
rect 3218 14660 3224 14662
rect 2916 14651 3224 14660
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2916 13628 3224 13637
rect 2916 13626 2922 13628
rect 2978 13626 3002 13628
rect 3058 13626 3082 13628
rect 3138 13626 3162 13628
rect 3218 13626 3224 13628
rect 2978 13574 2980 13626
rect 3160 13574 3162 13626
rect 2916 13572 2922 13574
rect 2978 13572 3002 13574
rect 3058 13572 3082 13574
rect 3138 13572 3162 13574
rect 3218 13572 3224 13574
rect 2916 13563 3224 13572
rect 3252 13258 3280 15302
rect 3608 15088 3660 15094
rect 3608 15030 3660 15036
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2608 12238 2636 12854
rect 2916 12540 3224 12549
rect 2916 12538 2922 12540
rect 2978 12538 3002 12540
rect 3058 12538 3082 12540
rect 3138 12538 3162 12540
rect 3218 12538 3224 12540
rect 2978 12486 2980 12538
rect 3160 12486 3162 12538
rect 2916 12484 2922 12486
rect 2978 12484 3002 12486
rect 3058 12484 3082 12486
rect 3138 12484 3162 12486
rect 3218 12484 3224 12486
rect 2916 12475 3224 12484
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2240 10198 2268 10610
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 2240 9586 2268 10134
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2424 9450 2452 11086
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1872 8974 1900 9318
rect 2608 9178 2636 11630
rect 2916 11452 3224 11461
rect 2916 11450 2922 11452
rect 2978 11450 3002 11452
rect 3058 11450 3082 11452
rect 3138 11450 3162 11452
rect 3218 11450 3224 11452
rect 2978 11398 2980 11450
rect 3160 11398 3162 11450
rect 2916 11396 2922 11398
rect 2978 11396 3002 11398
rect 3058 11396 3082 11398
rect 3138 11396 3162 11398
rect 3218 11396 3224 11398
rect 2916 11387 3224 11396
rect 3344 11354 3372 14894
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3436 11898 3464 13806
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3436 11354 3464 11698
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 11150 3556 12038
rect 3620 11286 3648 15030
rect 3712 14278 3740 15370
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3712 12986 3740 13126
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3804 12434 3832 15574
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 4882 15260 5190 15269
rect 4882 15258 4888 15260
rect 4944 15258 4968 15260
rect 5024 15258 5048 15260
rect 5104 15258 5128 15260
rect 5184 15258 5190 15260
rect 4944 15206 4946 15258
rect 5126 15206 5128 15258
rect 4882 15204 4888 15206
rect 4944 15204 4968 15206
rect 5024 15204 5048 15206
rect 5104 15204 5128 15206
rect 5184 15204 5190 15206
rect 4882 15195 5190 15204
rect 5736 15065 5764 15438
rect 5722 15056 5778 15065
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5632 15020 5684 15026
rect 5722 14991 5778 15000
rect 5816 15020 5868 15026
rect 5632 14962 5684 14968
rect 5816 14962 5868 14968
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3896 13734 3924 14350
rect 4882 14172 5190 14181
rect 4882 14170 4888 14172
rect 4944 14170 4968 14172
rect 5024 14170 5048 14172
rect 5104 14170 5128 14172
rect 5184 14170 5190 14172
rect 4944 14118 4946 14170
rect 5126 14118 5128 14170
rect 4882 14116 4888 14118
rect 4944 14116 4968 14118
rect 5024 14116 5048 14118
rect 5104 14116 5128 14118
rect 5184 14116 5190 14118
rect 4882 14107 5190 14116
rect 4160 14000 4212 14006
rect 4066 13968 4122 13977
rect 4160 13942 4212 13948
rect 4066 13903 4122 13912
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3896 13326 3924 13670
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3896 12986 3924 13262
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3712 12406 3832 12434
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10810 2820 11018
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 3712 10538 3740 12406
rect 4080 12238 4108 13903
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4080 11762 4108 12174
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3896 10674 3924 11698
rect 4080 11558 4108 11698
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 2916 10364 3224 10373
rect 2916 10362 2922 10364
rect 2978 10362 3002 10364
rect 3058 10362 3082 10364
rect 3138 10362 3162 10364
rect 3218 10362 3224 10364
rect 2978 10310 2980 10362
rect 3160 10310 3162 10362
rect 2916 10308 2922 10310
rect 2978 10308 3002 10310
rect 3058 10308 3082 10310
rect 3138 10308 3162 10310
rect 3218 10308 3224 10310
rect 2916 10299 3224 10308
rect 3712 9382 3740 10474
rect 4080 10470 4108 11494
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4172 10266 4200 13942
rect 5460 13734 5488 14962
rect 5644 13977 5672 14962
rect 5828 14634 5856 14962
rect 5736 14618 5856 14634
rect 5736 14612 5868 14618
rect 5736 14606 5816 14612
rect 5736 14006 5764 14606
rect 5816 14554 5868 14560
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5724 14000 5776 14006
rect 5630 13968 5686 13977
rect 5540 13932 5592 13938
rect 5724 13942 5776 13948
rect 5630 13903 5632 13912
rect 5540 13874 5592 13880
rect 5684 13903 5686 13912
rect 5632 13874 5684 13880
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4264 11898 4292 13194
rect 4448 12434 4476 13466
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12850 4660 13330
rect 4882 13084 5190 13093
rect 4882 13082 4888 13084
rect 4944 13082 4968 13084
rect 5024 13082 5048 13084
rect 5104 13082 5128 13084
rect 5184 13082 5190 13084
rect 4944 13030 4946 13082
rect 5126 13030 5128 13082
rect 4882 13028 4888 13030
rect 4944 13028 4968 13030
rect 5024 13028 5048 13030
rect 5104 13028 5128 13030
rect 5184 13028 5190 13030
rect 4882 13019 5190 13028
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 5172 12844 5224 12850
rect 5276 12832 5304 13670
rect 5224 12804 5304 12832
rect 5172 12786 5224 12792
rect 4620 12436 4672 12442
rect 4448 12406 4620 12434
rect 4620 12378 4672 12384
rect 4816 12322 4844 12786
rect 5276 12434 5304 12804
rect 5276 12406 5396 12434
rect 4724 12294 4844 12322
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4724 11626 4752 12294
rect 5368 12238 5396 12406
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10266 4292 11086
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10266 4568 10610
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 2916 9276 3224 9285
rect 2916 9274 2922 9276
rect 2978 9274 3002 9276
rect 3058 9274 3082 9276
rect 3138 9274 3162 9276
rect 3218 9274 3224 9276
rect 2978 9222 2980 9274
rect 3160 9222 3162 9274
rect 2916 9220 2922 9222
rect 2978 9220 3002 9222
rect 3058 9220 3082 9222
rect 3138 9220 3162 9222
rect 3218 9220 3224 9222
rect 2916 9211 3224 9220
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 2916 8188 3224 8197
rect 2916 8186 2922 8188
rect 2978 8186 3002 8188
rect 3058 8186 3082 8188
rect 3138 8186 3162 8188
rect 3218 8186 3224 8188
rect 2978 8134 2980 8186
rect 3160 8134 3162 8186
rect 2916 8132 2922 8134
rect 2978 8132 3002 8134
rect 3058 8132 3082 8134
rect 3138 8132 3162 8134
rect 3218 8132 3224 8134
rect 2916 8123 3224 8132
rect 2916 7100 3224 7109
rect 2916 7098 2922 7100
rect 2978 7098 3002 7100
rect 3058 7098 3082 7100
rect 3138 7098 3162 7100
rect 3218 7098 3224 7100
rect 2978 7046 2980 7098
rect 3160 7046 3162 7098
rect 2916 7044 2922 7046
rect 2978 7044 3002 7046
rect 3058 7044 3082 7046
rect 3138 7044 3162 7046
rect 3218 7044 3224 7046
rect 2916 7035 3224 7044
rect 4264 6730 4292 10202
rect 4724 9994 4752 11562
rect 4816 10810 4844 12174
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 4882 11996 5190 12005
rect 4882 11994 4888 11996
rect 4944 11994 4968 11996
rect 5024 11994 5048 11996
rect 5104 11994 5128 11996
rect 5184 11994 5190 11996
rect 4944 11942 4946 11994
rect 5126 11942 5128 11994
rect 4882 11940 4888 11942
rect 4944 11940 4968 11942
rect 5024 11940 5048 11942
rect 5104 11940 5128 11942
rect 5184 11940 5190 11942
rect 4882 11931 5190 11940
rect 5276 11898 5304 12038
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5368 11830 5396 12174
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5460 11762 5488 13670
rect 5552 12986 5580 13874
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12306 5672 12786
rect 5736 12782 5764 13330
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5736 12306 5764 12718
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 4882 10908 5190 10917
rect 4882 10906 4888 10908
rect 4944 10906 4968 10908
rect 5024 10906 5048 10908
rect 5104 10906 5128 10908
rect 5184 10906 5190 10908
rect 4944 10854 4946 10906
rect 5126 10854 5128 10906
rect 4882 10852 4888 10854
rect 4944 10852 4968 10854
rect 5024 10852 5048 10854
rect 5104 10852 5128 10854
rect 5184 10852 5190 10854
rect 4882 10843 5190 10852
rect 5552 10810 5580 11766
rect 5828 11286 5856 14418
rect 6012 14006 6040 15438
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 15162 6592 15302
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6550 15056 6606 15065
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 6288 13530 6316 15030
rect 6550 14991 6552 15000
rect 6604 14991 6606 15000
rect 6552 14962 6604 14968
rect 6564 14414 6592 14962
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6564 13326 6592 14350
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6656 14006 6684 14214
rect 6748 14074 6776 15438
rect 6849 14716 7157 14725
rect 6849 14714 6855 14716
rect 6911 14714 6935 14716
rect 6991 14714 7015 14716
rect 7071 14714 7095 14716
rect 7151 14714 7157 14716
rect 6911 14662 6913 14714
rect 7093 14662 7095 14714
rect 6849 14660 6855 14662
rect 6911 14660 6935 14662
rect 6991 14660 7015 14662
rect 7071 14660 7095 14662
rect 7151 14660 7157 14662
rect 6849 14651 7157 14660
rect 7576 14618 7604 15438
rect 8312 15162 8340 15438
rect 8815 15260 9123 15269
rect 8815 15258 8821 15260
rect 8877 15258 8901 15260
rect 8957 15258 8981 15260
rect 9037 15258 9061 15260
rect 9117 15258 9123 15260
rect 8877 15206 8879 15258
rect 9059 15206 9061 15258
rect 8815 15204 8821 15206
rect 8877 15204 8901 15206
rect 8957 15204 8981 15206
rect 9037 15204 9061 15206
rect 9117 15204 9123 15206
rect 8815 15195 9123 15204
rect 12748 15260 13056 15269
rect 12748 15258 12754 15260
rect 12810 15258 12834 15260
rect 12890 15258 12914 15260
rect 12970 15258 12994 15260
rect 13050 15258 13056 15260
rect 12810 15206 12812 15258
rect 12992 15206 12994 15258
rect 12748 15204 12754 15206
rect 12810 15204 12834 15206
rect 12890 15204 12914 15206
rect 12970 15204 12994 15206
rect 13050 15204 13056 15206
rect 12748 15195 13056 15204
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 10782 14716 11090 14725
rect 10782 14714 10788 14716
rect 10844 14714 10868 14716
rect 10924 14714 10948 14716
rect 11004 14714 11028 14716
rect 11084 14714 11090 14716
rect 10844 14662 10846 14714
rect 11026 14662 11028 14714
rect 10782 14660 10788 14662
rect 10844 14660 10868 14662
rect 10924 14660 10948 14662
rect 11004 14660 11028 14662
rect 11084 14660 11090 14662
rect 10782 14651 11090 14660
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6656 13326 6684 13942
rect 6840 13818 6868 14554
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 6748 13790 6868 13818
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6196 12918 6224 13262
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6288 11830 6316 13262
rect 6656 12850 6684 13262
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12238 6408 12582
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6748 12102 6776 13790
rect 6849 13628 7157 13637
rect 6849 13626 6855 13628
rect 6911 13626 6935 13628
rect 6991 13626 7015 13628
rect 7071 13626 7095 13628
rect 7151 13626 7157 13628
rect 6911 13574 6913 13626
rect 7093 13574 7095 13626
rect 6849 13572 6855 13574
rect 6911 13572 6935 13574
rect 6991 13572 7015 13574
rect 7071 13572 7095 13574
rect 7151 13572 7157 13574
rect 6849 13563 7157 13572
rect 7208 13394 7236 13874
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7300 13530 7328 13806
rect 7760 13530 7788 14350
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 13977 7880 14214
rect 8815 14172 9123 14181
rect 8815 14170 8821 14172
rect 8877 14170 8901 14172
rect 8957 14170 8981 14172
rect 9037 14170 9061 14172
rect 9117 14170 9123 14172
rect 8877 14118 8879 14170
rect 9059 14118 9061 14170
rect 8815 14116 8821 14118
rect 8877 14116 8901 14118
rect 8957 14116 8981 14118
rect 9037 14116 9061 14118
rect 9117 14116 9123 14118
rect 8815 14107 9123 14116
rect 12748 14172 13056 14181
rect 12748 14170 12754 14172
rect 12810 14170 12834 14172
rect 12890 14170 12914 14172
rect 12970 14170 12994 14172
rect 13050 14170 13056 14172
rect 12810 14118 12812 14170
rect 12992 14118 12994 14170
rect 12748 14116 12754 14118
rect 12810 14116 12834 14118
rect 12890 14116 12914 14118
rect 12970 14116 12994 14118
rect 13050 14116 13056 14118
rect 12748 14107 13056 14116
rect 7838 13968 7894 13977
rect 7838 13903 7894 13912
rect 10782 13628 11090 13637
rect 10782 13626 10788 13628
rect 10844 13626 10868 13628
rect 10924 13626 10948 13628
rect 11004 13626 11028 13628
rect 11084 13626 11090 13628
rect 10844 13574 10846 13626
rect 11026 13574 11028 13626
rect 10782 13572 10788 13574
rect 10844 13572 10868 13574
rect 10924 13572 10948 13574
rect 11004 13572 11028 13574
rect 11084 13572 11090 13574
rect 10782 13563 11090 13572
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7208 12646 7236 13330
rect 7300 12850 7328 13466
rect 8815 13084 9123 13093
rect 8815 13082 8821 13084
rect 8877 13082 8901 13084
rect 8957 13082 8981 13084
rect 9037 13082 9061 13084
rect 9117 13082 9123 13084
rect 8877 13030 8879 13082
rect 9059 13030 9061 13082
rect 8815 13028 8821 13030
rect 8877 13028 8901 13030
rect 8957 13028 8981 13030
rect 9037 13028 9061 13030
rect 9117 13028 9123 13030
rect 8815 13019 9123 13028
rect 12748 13084 13056 13093
rect 12748 13082 12754 13084
rect 12810 13082 12834 13084
rect 12890 13082 12914 13084
rect 12970 13082 12994 13084
rect 13050 13082 13056 13084
rect 12810 13030 12812 13082
rect 12992 13030 12994 13082
rect 12748 13028 12754 13030
rect 12810 13028 12834 13030
rect 12890 13028 12914 13030
rect 12970 13028 12994 13030
rect 13050 13028 13056 13030
rect 12748 13019 13056 13028
rect 7288 12844 7340 12850
rect 7340 12804 7420 12832
rect 7288 12786 7340 12792
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 6849 12540 7157 12549
rect 6849 12538 6855 12540
rect 6911 12538 6935 12540
rect 6991 12538 7015 12540
rect 7071 12538 7095 12540
rect 7151 12538 7157 12540
rect 6911 12486 6913 12538
rect 7093 12486 7095 12538
rect 6849 12484 6855 12486
rect 6911 12484 6935 12486
rect 6991 12484 7015 12486
rect 7071 12484 7095 12486
rect 7151 12484 7157 12486
rect 6849 12475 7157 12484
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5920 11286 5948 11630
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 6012 11218 6040 11494
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 10810 5672 11086
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 6012 10742 6040 11154
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6748 10674 6776 12038
rect 6849 11452 7157 11461
rect 6849 11450 6855 11452
rect 6911 11450 6935 11452
rect 6991 11450 7015 11452
rect 7071 11450 7095 11452
rect 7151 11450 7157 11452
rect 6911 11398 6913 11450
rect 7093 11398 7095 11450
rect 6849 11396 6855 11398
rect 6911 11396 6935 11398
rect 6991 11396 7015 11398
rect 7071 11396 7095 11398
rect 7151 11396 7157 11398
rect 6849 11387 7157 11396
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6748 10198 6776 10610
rect 6849 10364 7157 10373
rect 6849 10362 6855 10364
rect 6911 10362 6935 10364
rect 6991 10362 7015 10364
rect 7071 10362 7095 10364
rect 7151 10362 7157 10364
rect 6911 10310 6913 10362
rect 7093 10310 7095 10362
rect 6849 10308 6855 10310
rect 6911 10308 6935 10310
rect 6991 10308 7015 10310
rect 7071 10308 7095 10310
rect 7151 10308 7157 10310
rect 6849 10299 7157 10308
rect 7208 10266 7236 11018
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 7392 10130 7420 12804
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7484 10062 7512 12718
rect 10782 12540 11090 12549
rect 10782 12538 10788 12540
rect 10844 12538 10868 12540
rect 10924 12538 10948 12540
rect 11004 12538 11028 12540
rect 11084 12538 11090 12540
rect 10844 12486 10846 12538
rect 11026 12486 11028 12538
rect 10782 12484 10788 12486
rect 10844 12484 10868 12486
rect 10924 12484 10948 12486
rect 11004 12484 11028 12486
rect 11084 12484 11090 12486
rect 10782 12475 11090 12484
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8588 11762 8616 12038
rect 8815 11996 9123 12005
rect 8815 11994 8821 11996
rect 8877 11994 8901 11996
rect 8957 11994 8981 11996
rect 9037 11994 9061 11996
rect 9117 11994 9123 11996
rect 8877 11942 8879 11994
rect 9059 11942 9061 11994
rect 8815 11940 8821 11942
rect 8877 11940 8901 11942
rect 8957 11940 8981 11942
rect 9037 11940 9061 11942
rect 9117 11940 9123 11942
rect 8815 11931 9123 11940
rect 12748 11996 13056 12005
rect 12748 11994 12754 11996
rect 12810 11994 12834 11996
rect 12890 11994 12914 11996
rect 12970 11994 12994 11996
rect 13050 11994 13056 11996
rect 12810 11942 12812 11994
rect 12992 11942 12994 11994
rect 12748 11940 12754 11942
rect 12810 11940 12834 11942
rect 12890 11940 12914 11942
rect 12970 11940 12994 11942
rect 13050 11940 13056 11942
rect 12748 11931 13056 11940
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 8815 10908 9123 10917
rect 8815 10906 8821 10908
rect 8877 10906 8901 10908
rect 8957 10906 8981 10908
rect 9037 10906 9061 10908
rect 9117 10906 9123 10908
rect 8877 10854 8879 10906
rect 9059 10854 9061 10906
rect 8815 10852 8821 10854
rect 8877 10852 8901 10854
rect 8957 10852 8981 10854
rect 9037 10852 9061 10854
rect 9117 10852 9123 10854
rect 8815 10843 9123 10852
rect 9600 10606 9628 11494
rect 10782 11452 11090 11461
rect 10782 11450 10788 11452
rect 10844 11450 10868 11452
rect 10924 11450 10948 11452
rect 11004 11450 11028 11452
rect 11084 11450 11090 11452
rect 10844 11398 10846 11450
rect 11026 11398 11028 11450
rect 10782 11396 10788 11398
rect 10844 11396 10868 11398
rect 10924 11396 10948 11398
rect 11004 11396 11028 11398
rect 11084 11396 11090 11398
rect 10782 11387 11090 11396
rect 13372 11354 13400 17200
rect 14715 15804 15023 15813
rect 14715 15802 14721 15804
rect 14777 15802 14801 15804
rect 14857 15802 14881 15804
rect 14937 15802 14961 15804
rect 15017 15802 15023 15804
rect 14777 15750 14779 15802
rect 14959 15750 14961 15802
rect 14715 15748 14721 15750
rect 14777 15748 14801 15750
rect 14857 15748 14881 15750
rect 14937 15748 14961 15750
rect 15017 15748 15023 15750
rect 14715 15739 15023 15748
rect 16224 15706 16252 17326
rect 16302 17200 16358 17326
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16681 15260 16989 15269
rect 16681 15258 16687 15260
rect 16743 15258 16767 15260
rect 16823 15258 16847 15260
rect 16903 15258 16927 15260
rect 16983 15258 16989 15260
rect 16743 15206 16745 15258
rect 16925 15206 16927 15258
rect 16681 15204 16687 15206
rect 16743 15204 16767 15206
rect 16823 15204 16847 15206
rect 16903 15204 16927 15206
rect 16983 15204 16989 15206
rect 16681 15195 16989 15204
rect 14715 14716 15023 14725
rect 14715 14714 14721 14716
rect 14777 14714 14801 14716
rect 14857 14714 14881 14716
rect 14937 14714 14961 14716
rect 15017 14714 15023 14716
rect 14777 14662 14779 14714
rect 14959 14662 14961 14714
rect 14715 14660 14721 14662
rect 14777 14660 14801 14662
rect 14857 14660 14881 14662
rect 14937 14660 14961 14662
rect 15017 14660 15023 14662
rect 14715 14651 15023 14660
rect 16681 14172 16989 14181
rect 16681 14170 16687 14172
rect 16743 14170 16767 14172
rect 16823 14170 16847 14172
rect 16903 14170 16927 14172
rect 16983 14170 16989 14172
rect 16743 14118 16745 14170
rect 16925 14118 16927 14170
rect 16681 14116 16687 14118
rect 16743 14116 16767 14118
rect 16823 14116 16847 14118
rect 16903 14116 16927 14118
rect 16983 14116 16989 14118
rect 16681 14107 16989 14116
rect 14715 13628 15023 13637
rect 14715 13626 14721 13628
rect 14777 13626 14801 13628
rect 14857 13626 14881 13628
rect 14937 13626 14961 13628
rect 15017 13626 15023 13628
rect 14777 13574 14779 13626
rect 14959 13574 14961 13626
rect 14715 13572 14721 13574
rect 14777 13572 14801 13574
rect 14857 13572 14881 13574
rect 14937 13572 14961 13574
rect 15017 13572 15023 13574
rect 14715 13563 15023 13572
rect 16681 13084 16989 13093
rect 16681 13082 16687 13084
rect 16743 13082 16767 13084
rect 16823 13082 16847 13084
rect 16903 13082 16927 13084
rect 16983 13082 16989 13084
rect 16743 13030 16745 13082
rect 16925 13030 16927 13082
rect 16681 13028 16687 13030
rect 16743 13028 16767 13030
rect 16823 13028 16847 13030
rect 16903 13028 16927 13030
rect 16983 13028 16989 13030
rect 16681 13019 16989 13028
rect 14715 12540 15023 12549
rect 14715 12538 14721 12540
rect 14777 12538 14801 12540
rect 14857 12538 14881 12540
rect 14937 12538 14961 12540
rect 15017 12538 15023 12540
rect 14777 12486 14779 12538
rect 14959 12486 14961 12538
rect 14715 12484 14721 12486
rect 14777 12484 14801 12486
rect 14857 12484 14881 12486
rect 14937 12484 14961 12486
rect 15017 12484 15023 12486
rect 14715 12475 15023 12484
rect 16681 11996 16989 12005
rect 16681 11994 16687 11996
rect 16743 11994 16767 11996
rect 16823 11994 16847 11996
rect 16903 11994 16927 11996
rect 16983 11994 16989 11996
rect 16743 11942 16745 11994
rect 16925 11942 16927 11994
rect 16681 11940 16687 11942
rect 16743 11940 16767 11942
rect 16823 11940 16847 11942
rect 16903 11940 16927 11942
rect 16983 11940 16989 11942
rect 16681 11931 16989 11940
rect 14715 11452 15023 11461
rect 14715 11450 14721 11452
rect 14777 11450 14801 11452
rect 14857 11450 14881 11452
rect 14937 11450 14961 11452
rect 15017 11450 15023 11452
rect 14777 11398 14779 11450
rect 14959 11398 14961 11450
rect 14715 11396 14721 11398
rect 14777 11396 14801 11398
rect 14857 11396 14881 11398
rect 14937 11396 14961 11398
rect 15017 11396 15023 11398
rect 14715 11387 15023 11396
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 12748 10908 13056 10917
rect 12748 10906 12754 10908
rect 12810 10906 12834 10908
rect 12890 10906 12914 10908
rect 12970 10906 12994 10908
rect 13050 10906 13056 10908
rect 12810 10854 12812 10906
rect 12992 10854 12994 10906
rect 12748 10852 12754 10854
rect 12810 10852 12834 10854
rect 12890 10852 12914 10854
rect 12970 10852 12994 10854
rect 13050 10852 13056 10854
rect 12748 10843 13056 10852
rect 16681 10908 16989 10917
rect 16681 10906 16687 10908
rect 16743 10906 16767 10908
rect 16823 10906 16847 10908
rect 16903 10906 16927 10908
rect 16983 10906 16989 10908
rect 16743 10854 16745 10906
rect 16925 10854 16927 10906
rect 16681 10852 16687 10854
rect 16743 10852 16767 10854
rect 16823 10852 16847 10854
rect 16903 10852 16927 10854
rect 16983 10852 16989 10854
rect 16681 10843 16989 10852
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 10782 10364 11090 10373
rect 10782 10362 10788 10364
rect 10844 10362 10868 10364
rect 10924 10362 10948 10364
rect 11004 10362 11028 10364
rect 11084 10362 11090 10364
rect 10844 10310 10846 10362
rect 11026 10310 11028 10362
rect 10782 10308 10788 10310
rect 10844 10308 10868 10310
rect 10924 10308 10948 10310
rect 11004 10308 11028 10310
rect 11084 10308 11090 10310
rect 10782 10299 11090 10308
rect 14715 10364 15023 10373
rect 14715 10362 14721 10364
rect 14777 10362 14801 10364
rect 14857 10362 14881 10364
rect 14937 10362 14961 10364
rect 15017 10362 15023 10364
rect 14777 10310 14779 10362
rect 14959 10310 14961 10362
rect 14715 10308 14721 10310
rect 14777 10308 14801 10310
rect 14857 10308 14881 10310
rect 14937 10308 14961 10310
rect 15017 10308 15023 10310
rect 14715 10299 15023 10308
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4724 9518 4752 9930
rect 4882 9820 5190 9829
rect 4882 9818 4888 9820
rect 4944 9818 4968 9820
rect 5024 9818 5048 9820
rect 5104 9818 5128 9820
rect 5184 9818 5190 9820
rect 4944 9766 4946 9818
rect 5126 9766 5128 9818
rect 4882 9764 4888 9766
rect 4944 9764 4968 9766
rect 5024 9764 5048 9766
rect 5104 9764 5128 9766
rect 5184 9764 5190 9766
rect 4882 9755 5190 9764
rect 8815 9820 9123 9829
rect 8815 9818 8821 9820
rect 8877 9818 8901 9820
rect 8957 9818 8981 9820
rect 9037 9818 9061 9820
rect 9117 9818 9123 9820
rect 8877 9766 8879 9818
rect 9059 9766 9061 9818
rect 8815 9764 8821 9766
rect 8877 9764 8901 9766
rect 8957 9764 8981 9766
rect 9037 9764 9061 9766
rect 9117 9764 9123 9766
rect 8815 9755 9123 9764
rect 12748 9820 13056 9829
rect 12748 9818 12754 9820
rect 12810 9818 12834 9820
rect 12890 9818 12914 9820
rect 12970 9818 12994 9820
rect 13050 9818 13056 9820
rect 12810 9766 12812 9818
rect 12992 9766 12994 9818
rect 12748 9764 12754 9766
rect 12810 9764 12834 9766
rect 12890 9764 12914 9766
rect 12970 9764 12994 9766
rect 13050 9764 13056 9766
rect 12748 9755 13056 9764
rect 16681 9820 16989 9829
rect 16681 9818 16687 9820
rect 16743 9818 16767 9820
rect 16823 9818 16847 9820
rect 16903 9818 16927 9820
rect 16983 9818 16989 9820
rect 16743 9766 16745 9818
rect 16925 9766 16927 9818
rect 16681 9764 16687 9766
rect 16743 9764 16767 9766
rect 16823 9764 16847 9766
rect 16903 9764 16927 9766
rect 16983 9764 16989 9766
rect 16681 9755 16989 9764
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 6849 9276 7157 9285
rect 6849 9274 6855 9276
rect 6911 9274 6935 9276
rect 6991 9274 7015 9276
rect 7071 9274 7095 9276
rect 7151 9274 7157 9276
rect 6911 9222 6913 9274
rect 7093 9222 7095 9274
rect 6849 9220 6855 9222
rect 6911 9220 6935 9222
rect 6991 9220 7015 9222
rect 7071 9220 7095 9222
rect 7151 9220 7157 9222
rect 6849 9211 7157 9220
rect 10782 9276 11090 9285
rect 10782 9274 10788 9276
rect 10844 9274 10868 9276
rect 10924 9274 10948 9276
rect 11004 9274 11028 9276
rect 11084 9274 11090 9276
rect 10844 9222 10846 9274
rect 11026 9222 11028 9274
rect 10782 9220 10788 9222
rect 10844 9220 10868 9222
rect 10924 9220 10948 9222
rect 11004 9220 11028 9222
rect 11084 9220 11090 9222
rect 10782 9211 11090 9220
rect 14715 9276 15023 9285
rect 14715 9274 14721 9276
rect 14777 9274 14801 9276
rect 14857 9274 14881 9276
rect 14937 9274 14961 9276
rect 15017 9274 15023 9276
rect 14777 9222 14779 9274
rect 14959 9222 14961 9274
rect 14715 9220 14721 9222
rect 14777 9220 14801 9222
rect 14857 9220 14881 9222
rect 14937 9220 14961 9222
rect 15017 9220 15023 9222
rect 14715 9211 15023 9220
rect 4882 8732 5190 8741
rect 4882 8730 4888 8732
rect 4944 8730 4968 8732
rect 5024 8730 5048 8732
rect 5104 8730 5128 8732
rect 5184 8730 5190 8732
rect 4944 8678 4946 8730
rect 5126 8678 5128 8730
rect 4882 8676 4888 8678
rect 4944 8676 4968 8678
rect 5024 8676 5048 8678
rect 5104 8676 5128 8678
rect 5184 8676 5190 8678
rect 4882 8667 5190 8676
rect 8815 8732 9123 8741
rect 8815 8730 8821 8732
rect 8877 8730 8901 8732
rect 8957 8730 8981 8732
rect 9037 8730 9061 8732
rect 9117 8730 9123 8732
rect 8877 8678 8879 8730
rect 9059 8678 9061 8730
rect 8815 8676 8821 8678
rect 8877 8676 8901 8678
rect 8957 8676 8981 8678
rect 9037 8676 9061 8678
rect 9117 8676 9123 8678
rect 8815 8667 9123 8676
rect 12748 8732 13056 8741
rect 12748 8730 12754 8732
rect 12810 8730 12834 8732
rect 12890 8730 12914 8732
rect 12970 8730 12994 8732
rect 13050 8730 13056 8732
rect 12810 8678 12812 8730
rect 12992 8678 12994 8730
rect 12748 8676 12754 8678
rect 12810 8676 12834 8678
rect 12890 8676 12914 8678
rect 12970 8676 12994 8678
rect 13050 8676 13056 8678
rect 12748 8667 13056 8676
rect 16681 8732 16989 8741
rect 16681 8730 16687 8732
rect 16743 8730 16767 8732
rect 16823 8730 16847 8732
rect 16903 8730 16927 8732
rect 16983 8730 16989 8732
rect 16743 8678 16745 8730
rect 16925 8678 16927 8730
rect 16681 8676 16687 8678
rect 16743 8676 16767 8678
rect 16823 8676 16847 8678
rect 16903 8676 16927 8678
rect 16983 8676 16989 8678
rect 16681 8667 16989 8676
rect 6849 8188 7157 8197
rect 6849 8186 6855 8188
rect 6911 8186 6935 8188
rect 6991 8186 7015 8188
rect 7071 8186 7095 8188
rect 7151 8186 7157 8188
rect 6911 8134 6913 8186
rect 7093 8134 7095 8186
rect 6849 8132 6855 8134
rect 6911 8132 6935 8134
rect 6991 8132 7015 8134
rect 7071 8132 7095 8134
rect 7151 8132 7157 8134
rect 6849 8123 7157 8132
rect 10782 8188 11090 8197
rect 10782 8186 10788 8188
rect 10844 8186 10868 8188
rect 10924 8186 10948 8188
rect 11004 8186 11028 8188
rect 11084 8186 11090 8188
rect 10844 8134 10846 8186
rect 11026 8134 11028 8186
rect 10782 8132 10788 8134
rect 10844 8132 10868 8134
rect 10924 8132 10948 8134
rect 11004 8132 11028 8134
rect 11084 8132 11090 8134
rect 10782 8123 11090 8132
rect 14715 8188 15023 8197
rect 14715 8186 14721 8188
rect 14777 8186 14801 8188
rect 14857 8186 14881 8188
rect 14937 8186 14961 8188
rect 15017 8186 15023 8188
rect 14777 8134 14779 8186
rect 14959 8134 14961 8186
rect 14715 8132 14721 8134
rect 14777 8132 14801 8134
rect 14857 8132 14881 8134
rect 14937 8132 14961 8134
rect 15017 8132 15023 8134
rect 14715 8123 15023 8132
rect 4882 7644 5190 7653
rect 4882 7642 4888 7644
rect 4944 7642 4968 7644
rect 5024 7642 5048 7644
rect 5104 7642 5128 7644
rect 5184 7642 5190 7644
rect 4944 7590 4946 7642
rect 5126 7590 5128 7642
rect 4882 7588 4888 7590
rect 4944 7588 4968 7590
rect 5024 7588 5048 7590
rect 5104 7588 5128 7590
rect 5184 7588 5190 7590
rect 4882 7579 5190 7588
rect 8815 7644 9123 7653
rect 8815 7642 8821 7644
rect 8877 7642 8901 7644
rect 8957 7642 8981 7644
rect 9037 7642 9061 7644
rect 9117 7642 9123 7644
rect 8877 7590 8879 7642
rect 9059 7590 9061 7642
rect 8815 7588 8821 7590
rect 8877 7588 8901 7590
rect 8957 7588 8981 7590
rect 9037 7588 9061 7590
rect 9117 7588 9123 7590
rect 8815 7579 9123 7588
rect 12748 7644 13056 7653
rect 12748 7642 12754 7644
rect 12810 7642 12834 7644
rect 12890 7642 12914 7644
rect 12970 7642 12994 7644
rect 13050 7642 13056 7644
rect 12810 7590 12812 7642
rect 12992 7590 12994 7642
rect 12748 7588 12754 7590
rect 12810 7588 12834 7590
rect 12890 7588 12914 7590
rect 12970 7588 12994 7590
rect 13050 7588 13056 7590
rect 12748 7579 13056 7588
rect 16681 7644 16989 7653
rect 16681 7642 16687 7644
rect 16743 7642 16767 7644
rect 16823 7642 16847 7644
rect 16903 7642 16927 7644
rect 16983 7642 16989 7644
rect 16743 7590 16745 7642
rect 16925 7590 16927 7642
rect 16681 7588 16687 7590
rect 16743 7588 16767 7590
rect 16823 7588 16847 7590
rect 16903 7588 16927 7590
rect 16983 7588 16989 7590
rect 16681 7579 16989 7588
rect 6849 7100 7157 7109
rect 6849 7098 6855 7100
rect 6911 7098 6935 7100
rect 6991 7098 7015 7100
rect 7071 7098 7095 7100
rect 7151 7098 7157 7100
rect 6911 7046 6913 7098
rect 7093 7046 7095 7098
rect 6849 7044 6855 7046
rect 6911 7044 6935 7046
rect 6991 7044 7015 7046
rect 7071 7044 7095 7046
rect 7151 7044 7157 7046
rect 6849 7035 7157 7044
rect 10782 7100 11090 7109
rect 10782 7098 10788 7100
rect 10844 7098 10868 7100
rect 10924 7098 10948 7100
rect 11004 7098 11028 7100
rect 11084 7098 11090 7100
rect 10844 7046 10846 7098
rect 11026 7046 11028 7098
rect 10782 7044 10788 7046
rect 10844 7044 10868 7046
rect 10924 7044 10948 7046
rect 11004 7044 11028 7046
rect 11084 7044 11090 7046
rect 10782 7035 11090 7044
rect 14715 7100 15023 7109
rect 14715 7098 14721 7100
rect 14777 7098 14801 7100
rect 14857 7098 14881 7100
rect 14937 7098 14961 7100
rect 15017 7098 15023 7100
rect 14777 7046 14779 7098
rect 14959 7046 14961 7098
rect 14715 7044 14721 7046
rect 14777 7044 14801 7046
rect 14857 7044 14881 7046
rect 14937 7044 14961 7046
rect 15017 7044 15023 7046
rect 14715 7035 15023 7044
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4882 6556 5190 6565
rect 4882 6554 4888 6556
rect 4944 6554 4968 6556
rect 5024 6554 5048 6556
rect 5104 6554 5128 6556
rect 5184 6554 5190 6556
rect 4944 6502 4946 6554
rect 5126 6502 5128 6554
rect 4882 6500 4888 6502
rect 4944 6500 4968 6502
rect 5024 6500 5048 6502
rect 5104 6500 5128 6502
rect 5184 6500 5190 6502
rect 4882 6491 5190 6500
rect 8815 6556 9123 6565
rect 8815 6554 8821 6556
rect 8877 6554 8901 6556
rect 8957 6554 8981 6556
rect 9037 6554 9061 6556
rect 9117 6554 9123 6556
rect 8877 6502 8879 6554
rect 9059 6502 9061 6554
rect 8815 6500 8821 6502
rect 8877 6500 8901 6502
rect 8957 6500 8981 6502
rect 9037 6500 9061 6502
rect 9117 6500 9123 6502
rect 8815 6491 9123 6500
rect 12748 6556 13056 6565
rect 12748 6554 12754 6556
rect 12810 6554 12834 6556
rect 12890 6554 12914 6556
rect 12970 6554 12994 6556
rect 13050 6554 13056 6556
rect 12810 6502 12812 6554
rect 12992 6502 12994 6554
rect 12748 6500 12754 6502
rect 12810 6500 12834 6502
rect 12890 6500 12914 6502
rect 12970 6500 12994 6502
rect 13050 6500 13056 6502
rect 12748 6491 13056 6500
rect 16681 6556 16989 6565
rect 16681 6554 16687 6556
rect 16743 6554 16767 6556
rect 16823 6554 16847 6556
rect 16903 6554 16927 6556
rect 16983 6554 16989 6556
rect 16743 6502 16745 6554
rect 16925 6502 16927 6554
rect 16681 6500 16687 6502
rect 16743 6500 16767 6502
rect 16823 6500 16847 6502
rect 16903 6500 16927 6502
rect 16983 6500 16989 6502
rect 16681 6491 16989 6500
rect 2916 6012 3224 6021
rect 2916 6010 2922 6012
rect 2978 6010 3002 6012
rect 3058 6010 3082 6012
rect 3138 6010 3162 6012
rect 3218 6010 3224 6012
rect 2978 5958 2980 6010
rect 3160 5958 3162 6010
rect 2916 5956 2922 5958
rect 2978 5956 3002 5958
rect 3058 5956 3082 5958
rect 3138 5956 3162 5958
rect 3218 5956 3224 5958
rect 2916 5947 3224 5956
rect 6849 6012 7157 6021
rect 6849 6010 6855 6012
rect 6911 6010 6935 6012
rect 6991 6010 7015 6012
rect 7071 6010 7095 6012
rect 7151 6010 7157 6012
rect 6911 5958 6913 6010
rect 7093 5958 7095 6010
rect 6849 5956 6855 5958
rect 6911 5956 6935 5958
rect 6991 5956 7015 5958
rect 7071 5956 7095 5958
rect 7151 5956 7157 5958
rect 6849 5947 7157 5956
rect 10782 6012 11090 6021
rect 10782 6010 10788 6012
rect 10844 6010 10868 6012
rect 10924 6010 10948 6012
rect 11004 6010 11028 6012
rect 11084 6010 11090 6012
rect 10844 5958 10846 6010
rect 11026 5958 11028 6010
rect 10782 5956 10788 5958
rect 10844 5956 10868 5958
rect 10924 5956 10948 5958
rect 11004 5956 11028 5958
rect 11084 5956 11090 5958
rect 10782 5947 11090 5956
rect 14715 6012 15023 6021
rect 14715 6010 14721 6012
rect 14777 6010 14801 6012
rect 14857 6010 14881 6012
rect 14937 6010 14961 6012
rect 15017 6010 15023 6012
rect 14777 5958 14779 6010
rect 14959 5958 14961 6010
rect 14715 5956 14721 5958
rect 14777 5956 14801 5958
rect 14857 5956 14881 5958
rect 14937 5956 14961 5958
rect 15017 5956 15023 5958
rect 14715 5947 15023 5956
rect 4882 5468 5190 5477
rect 4882 5466 4888 5468
rect 4944 5466 4968 5468
rect 5024 5466 5048 5468
rect 5104 5466 5128 5468
rect 5184 5466 5190 5468
rect 4944 5414 4946 5466
rect 5126 5414 5128 5466
rect 4882 5412 4888 5414
rect 4944 5412 4968 5414
rect 5024 5412 5048 5414
rect 5104 5412 5128 5414
rect 5184 5412 5190 5414
rect 4882 5403 5190 5412
rect 8815 5468 9123 5477
rect 8815 5466 8821 5468
rect 8877 5466 8901 5468
rect 8957 5466 8981 5468
rect 9037 5466 9061 5468
rect 9117 5466 9123 5468
rect 8877 5414 8879 5466
rect 9059 5414 9061 5466
rect 8815 5412 8821 5414
rect 8877 5412 8901 5414
rect 8957 5412 8981 5414
rect 9037 5412 9061 5414
rect 9117 5412 9123 5414
rect 8815 5403 9123 5412
rect 12748 5468 13056 5477
rect 12748 5466 12754 5468
rect 12810 5466 12834 5468
rect 12890 5466 12914 5468
rect 12970 5466 12994 5468
rect 13050 5466 13056 5468
rect 12810 5414 12812 5466
rect 12992 5414 12994 5466
rect 12748 5412 12754 5414
rect 12810 5412 12834 5414
rect 12890 5412 12914 5414
rect 12970 5412 12994 5414
rect 13050 5412 13056 5414
rect 12748 5403 13056 5412
rect 16681 5468 16989 5477
rect 16681 5466 16687 5468
rect 16743 5466 16767 5468
rect 16823 5466 16847 5468
rect 16903 5466 16927 5468
rect 16983 5466 16989 5468
rect 16743 5414 16745 5466
rect 16925 5414 16927 5466
rect 16681 5412 16687 5414
rect 16743 5412 16767 5414
rect 16823 5412 16847 5414
rect 16903 5412 16927 5414
rect 16983 5412 16989 5414
rect 16681 5403 16989 5412
rect 2916 4924 3224 4933
rect 2916 4922 2922 4924
rect 2978 4922 3002 4924
rect 3058 4922 3082 4924
rect 3138 4922 3162 4924
rect 3218 4922 3224 4924
rect 2978 4870 2980 4922
rect 3160 4870 3162 4922
rect 2916 4868 2922 4870
rect 2978 4868 3002 4870
rect 3058 4868 3082 4870
rect 3138 4868 3162 4870
rect 3218 4868 3224 4870
rect 2916 4859 3224 4868
rect 6849 4924 7157 4933
rect 6849 4922 6855 4924
rect 6911 4922 6935 4924
rect 6991 4922 7015 4924
rect 7071 4922 7095 4924
rect 7151 4922 7157 4924
rect 6911 4870 6913 4922
rect 7093 4870 7095 4922
rect 6849 4868 6855 4870
rect 6911 4868 6935 4870
rect 6991 4868 7015 4870
rect 7071 4868 7095 4870
rect 7151 4868 7157 4870
rect 6849 4859 7157 4868
rect 10782 4924 11090 4933
rect 10782 4922 10788 4924
rect 10844 4922 10868 4924
rect 10924 4922 10948 4924
rect 11004 4922 11028 4924
rect 11084 4922 11090 4924
rect 10844 4870 10846 4922
rect 11026 4870 11028 4922
rect 10782 4868 10788 4870
rect 10844 4868 10868 4870
rect 10924 4868 10948 4870
rect 11004 4868 11028 4870
rect 11084 4868 11090 4870
rect 10782 4859 11090 4868
rect 14715 4924 15023 4933
rect 14715 4922 14721 4924
rect 14777 4922 14801 4924
rect 14857 4922 14881 4924
rect 14937 4922 14961 4924
rect 15017 4922 15023 4924
rect 14777 4870 14779 4922
rect 14959 4870 14961 4922
rect 14715 4868 14721 4870
rect 14777 4868 14801 4870
rect 14857 4868 14881 4870
rect 14937 4868 14961 4870
rect 15017 4868 15023 4870
rect 14715 4859 15023 4868
rect 4882 4380 5190 4389
rect 4882 4378 4888 4380
rect 4944 4378 4968 4380
rect 5024 4378 5048 4380
rect 5104 4378 5128 4380
rect 5184 4378 5190 4380
rect 4944 4326 4946 4378
rect 5126 4326 5128 4378
rect 4882 4324 4888 4326
rect 4944 4324 4968 4326
rect 5024 4324 5048 4326
rect 5104 4324 5128 4326
rect 5184 4324 5190 4326
rect 4882 4315 5190 4324
rect 8815 4380 9123 4389
rect 8815 4378 8821 4380
rect 8877 4378 8901 4380
rect 8957 4378 8981 4380
rect 9037 4378 9061 4380
rect 9117 4378 9123 4380
rect 8877 4326 8879 4378
rect 9059 4326 9061 4378
rect 8815 4324 8821 4326
rect 8877 4324 8901 4326
rect 8957 4324 8981 4326
rect 9037 4324 9061 4326
rect 9117 4324 9123 4326
rect 8815 4315 9123 4324
rect 12748 4380 13056 4389
rect 12748 4378 12754 4380
rect 12810 4378 12834 4380
rect 12890 4378 12914 4380
rect 12970 4378 12994 4380
rect 13050 4378 13056 4380
rect 12810 4326 12812 4378
rect 12992 4326 12994 4378
rect 12748 4324 12754 4326
rect 12810 4324 12834 4326
rect 12890 4324 12914 4326
rect 12970 4324 12994 4326
rect 13050 4324 13056 4326
rect 12748 4315 13056 4324
rect 16681 4380 16989 4389
rect 16681 4378 16687 4380
rect 16743 4378 16767 4380
rect 16823 4378 16847 4380
rect 16903 4378 16927 4380
rect 16983 4378 16989 4380
rect 16743 4326 16745 4378
rect 16925 4326 16927 4378
rect 16681 4324 16687 4326
rect 16743 4324 16767 4326
rect 16823 4324 16847 4326
rect 16903 4324 16927 4326
rect 16983 4324 16989 4326
rect 16681 4315 16989 4324
rect 2916 3836 3224 3845
rect 2916 3834 2922 3836
rect 2978 3834 3002 3836
rect 3058 3834 3082 3836
rect 3138 3834 3162 3836
rect 3218 3834 3224 3836
rect 2978 3782 2980 3834
rect 3160 3782 3162 3834
rect 2916 3780 2922 3782
rect 2978 3780 3002 3782
rect 3058 3780 3082 3782
rect 3138 3780 3162 3782
rect 3218 3780 3224 3782
rect 2916 3771 3224 3780
rect 6849 3836 7157 3845
rect 6849 3834 6855 3836
rect 6911 3834 6935 3836
rect 6991 3834 7015 3836
rect 7071 3834 7095 3836
rect 7151 3834 7157 3836
rect 6911 3782 6913 3834
rect 7093 3782 7095 3834
rect 6849 3780 6855 3782
rect 6911 3780 6935 3782
rect 6991 3780 7015 3782
rect 7071 3780 7095 3782
rect 7151 3780 7157 3782
rect 6849 3771 7157 3780
rect 10782 3836 11090 3845
rect 10782 3834 10788 3836
rect 10844 3834 10868 3836
rect 10924 3834 10948 3836
rect 11004 3834 11028 3836
rect 11084 3834 11090 3836
rect 10844 3782 10846 3834
rect 11026 3782 11028 3834
rect 10782 3780 10788 3782
rect 10844 3780 10868 3782
rect 10924 3780 10948 3782
rect 11004 3780 11028 3782
rect 11084 3780 11090 3782
rect 10782 3771 11090 3780
rect 14715 3836 15023 3845
rect 14715 3834 14721 3836
rect 14777 3834 14801 3836
rect 14857 3834 14881 3836
rect 14937 3834 14961 3836
rect 15017 3834 15023 3836
rect 14777 3782 14779 3834
rect 14959 3782 14961 3834
rect 14715 3780 14721 3782
rect 14777 3780 14801 3782
rect 14857 3780 14881 3782
rect 14937 3780 14961 3782
rect 15017 3780 15023 3782
rect 14715 3771 15023 3780
rect 4882 3292 5190 3301
rect 4882 3290 4888 3292
rect 4944 3290 4968 3292
rect 5024 3290 5048 3292
rect 5104 3290 5128 3292
rect 5184 3290 5190 3292
rect 4944 3238 4946 3290
rect 5126 3238 5128 3290
rect 4882 3236 4888 3238
rect 4944 3236 4968 3238
rect 5024 3236 5048 3238
rect 5104 3236 5128 3238
rect 5184 3236 5190 3238
rect 4882 3227 5190 3236
rect 8815 3292 9123 3301
rect 8815 3290 8821 3292
rect 8877 3290 8901 3292
rect 8957 3290 8981 3292
rect 9037 3290 9061 3292
rect 9117 3290 9123 3292
rect 8877 3238 8879 3290
rect 9059 3238 9061 3290
rect 8815 3236 8821 3238
rect 8877 3236 8901 3238
rect 8957 3236 8981 3238
rect 9037 3236 9061 3238
rect 9117 3236 9123 3238
rect 8815 3227 9123 3236
rect 12748 3292 13056 3301
rect 12748 3290 12754 3292
rect 12810 3290 12834 3292
rect 12890 3290 12914 3292
rect 12970 3290 12994 3292
rect 13050 3290 13056 3292
rect 12810 3238 12812 3290
rect 12992 3238 12994 3290
rect 12748 3236 12754 3238
rect 12810 3236 12834 3238
rect 12890 3236 12914 3238
rect 12970 3236 12994 3238
rect 13050 3236 13056 3238
rect 12748 3227 13056 3236
rect 16681 3292 16989 3301
rect 16681 3290 16687 3292
rect 16743 3290 16767 3292
rect 16823 3290 16847 3292
rect 16903 3290 16927 3292
rect 16983 3290 16989 3292
rect 16743 3238 16745 3290
rect 16925 3238 16927 3290
rect 16681 3236 16687 3238
rect 16743 3236 16767 3238
rect 16823 3236 16847 3238
rect 16903 3236 16927 3238
rect 16983 3236 16989 3238
rect 16681 3227 16989 3236
rect 2916 2748 3224 2757
rect 2916 2746 2922 2748
rect 2978 2746 3002 2748
rect 3058 2746 3082 2748
rect 3138 2746 3162 2748
rect 3218 2746 3224 2748
rect 2978 2694 2980 2746
rect 3160 2694 3162 2746
rect 2916 2692 2922 2694
rect 2978 2692 3002 2694
rect 3058 2692 3082 2694
rect 3138 2692 3162 2694
rect 3218 2692 3224 2694
rect 2916 2683 3224 2692
rect 6849 2748 7157 2757
rect 6849 2746 6855 2748
rect 6911 2746 6935 2748
rect 6991 2746 7015 2748
rect 7071 2746 7095 2748
rect 7151 2746 7157 2748
rect 6911 2694 6913 2746
rect 7093 2694 7095 2746
rect 6849 2692 6855 2694
rect 6911 2692 6935 2694
rect 6991 2692 7015 2694
rect 7071 2692 7095 2694
rect 7151 2692 7157 2694
rect 6849 2683 7157 2692
rect 10782 2748 11090 2757
rect 10782 2746 10788 2748
rect 10844 2746 10868 2748
rect 10924 2746 10948 2748
rect 11004 2746 11028 2748
rect 11084 2746 11090 2748
rect 10844 2694 10846 2746
rect 11026 2694 11028 2746
rect 10782 2692 10788 2694
rect 10844 2692 10868 2694
rect 10924 2692 10948 2694
rect 11004 2692 11028 2694
rect 11084 2692 11090 2694
rect 10782 2683 11090 2692
rect 14715 2748 15023 2757
rect 14715 2746 14721 2748
rect 14777 2746 14801 2748
rect 14857 2746 14881 2748
rect 14937 2746 14961 2748
rect 15017 2746 15023 2748
rect 14777 2694 14779 2746
rect 14959 2694 14961 2746
rect 14715 2692 14721 2694
rect 14777 2692 14801 2694
rect 14857 2692 14881 2694
rect 14937 2692 14961 2694
rect 15017 2692 15023 2694
rect 14715 2683 15023 2692
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1768 2304 1820 2310
rect 1766 2272 1768 2281
rect 1820 2272 1822 2281
rect 1766 2207 1822 2216
rect 4882 2204 5190 2213
rect 4882 2202 4888 2204
rect 4944 2202 4968 2204
rect 5024 2202 5048 2204
rect 5104 2202 5128 2204
rect 5184 2202 5190 2204
rect 4944 2150 4946 2202
rect 5126 2150 5128 2202
rect 4882 2148 4888 2150
rect 4944 2148 4968 2150
rect 5024 2148 5048 2150
rect 5104 2148 5128 2150
rect 5184 2148 5190 2150
rect 4882 2139 5190 2148
rect 8815 2204 9123 2213
rect 8815 2202 8821 2204
rect 8877 2202 8901 2204
rect 8957 2202 8981 2204
rect 9037 2202 9061 2204
rect 9117 2202 9123 2204
rect 8877 2150 8879 2202
rect 9059 2150 9061 2202
rect 8815 2148 8821 2150
rect 8877 2148 8901 2150
rect 8957 2148 8981 2150
rect 9037 2148 9061 2150
rect 9117 2148 9123 2150
rect 8815 2139 9123 2148
rect 12748 2204 13056 2213
rect 12748 2202 12754 2204
rect 12810 2202 12834 2204
rect 12890 2202 12914 2204
rect 12970 2202 12994 2204
rect 13050 2202 13056 2204
rect 12810 2150 12812 2202
rect 12992 2150 12994 2202
rect 12748 2148 12754 2150
rect 12810 2148 12834 2150
rect 12890 2148 12914 2150
rect 12970 2148 12994 2150
rect 13050 2148 13056 2150
rect 12748 2139 13056 2148
rect 16681 2204 16989 2213
rect 16681 2202 16687 2204
rect 16743 2202 16767 2204
rect 16823 2202 16847 2204
rect 16903 2202 16927 2204
rect 16983 2202 16989 2204
rect 16743 2150 16745 2202
rect 16925 2150 16927 2202
rect 16681 2148 16687 2150
rect 16743 2148 16767 2150
rect 16823 2148 16847 2150
rect 16903 2148 16927 2150
rect 16983 2148 16989 2150
rect 16681 2139 16989 2148
<< via2 >>
rect 2922 15802 2978 15804
rect 3002 15802 3058 15804
rect 3082 15802 3138 15804
rect 3162 15802 3218 15804
rect 2922 15750 2968 15802
rect 2968 15750 2978 15802
rect 3002 15750 3032 15802
rect 3032 15750 3044 15802
rect 3044 15750 3058 15802
rect 3082 15750 3096 15802
rect 3096 15750 3108 15802
rect 3108 15750 3138 15802
rect 3162 15750 3172 15802
rect 3172 15750 3218 15802
rect 2922 15748 2978 15750
rect 3002 15748 3058 15750
rect 3082 15748 3138 15750
rect 3162 15748 3218 15750
rect 2778 15680 2834 15736
rect 6855 15802 6911 15804
rect 6935 15802 6991 15804
rect 7015 15802 7071 15804
rect 7095 15802 7151 15804
rect 6855 15750 6901 15802
rect 6901 15750 6911 15802
rect 6935 15750 6965 15802
rect 6965 15750 6977 15802
rect 6977 15750 6991 15802
rect 7015 15750 7029 15802
rect 7029 15750 7041 15802
rect 7041 15750 7071 15802
rect 7095 15750 7105 15802
rect 7105 15750 7151 15802
rect 6855 15748 6911 15750
rect 6935 15748 6991 15750
rect 7015 15748 7071 15750
rect 7095 15748 7151 15750
rect 10788 15802 10844 15804
rect 10868 15802 10924 15804
rect 10948 15802 11004 15804
rect 11028 15802 11084 15804
rect 10788 15750 10834 15802
rect 10834 15750 10844 15802
rect 10868 15750 10898 15802
rect 10898 15750 10910 15802
rect 10910 15750 10924 15802
rect 10948 15750 10962 15802
rect 10962 15750 10974 15802
rect 10974 15750 11004 15802
rect 11028 15750 11038 15802
rect 11038 15750 11084 15802
rect 10788 15748 10844 15750
rect 10868 15748 10924 15750
rect 10948 15748 11004 15750
rect 11028 15748 11084 15750
rect 2226 13932 2282 13968
rect 2226 13912 2228 13932
rect 2228 13912 2280 13932
rect 2280 13912 2282 13932
rect 1490 6740 1492 6760
rect 1492 6740 1544 6760
rect 1544 6740 1546 6760
rect 1490 6704 1546 6740
rect 1674 11192 1730 11248
rect 2922 14714 2978 14716
rect 3002 14714 3058 14716
rect 3082 14714 3138 14716
rect 3162 14714 3218 14716
rect 2922 14662 2968 14714
rect 2968 14662 2978 14714
rect 3002 14662 3032 14714
rect 3032 14662 3044 14714
rect 3044 14662 3058 14714
rect 3082 14662 3096 14714
rect 3096 14662 3108 14714
rect 3108 14662 3138 14714
rect 3162 14662 3172 14714
rect 3172 14662 3218 14714
rect 2922 14660 2978 14662
rect 3002 14660 3058 14662
rect 3082 14660 3138 14662
rect 3162 14660 3218 14662
rect 2922 13626 2978 13628
rect 3002 13626 3058 13628
rect 3082 13626 3138 13628
rect 3162 13626 3218 13628
rect 2922 13574 2968 13626
rect 2968 13574 2978 13626
rect 3002 13574 3032 13626
rect 3032 13574 3044 13626
rect 3044 13574 3058 13626
rect 3082 13574 3096 13626
rect 3096 13574 3108 13626
rect 3108 13574 3138 13626
rect 3162 13574 3172 13626
rect 3172 13574 3218 13626
rect 2922 13572 2978 13574
rect 3002 13572 3058 13574
rect 3082 13572 3138 13574
rect 3162 13572 3218 13574
rect 2922 12538 2978 12540
rect 3002 12538 3058 12540
rect 3082 12538 3138 12540
rect 3162 12538 3218 12540
rect 2922 12486 2968 12538
rect 2968 12486 2978 12538
rect 3002 12486 3032 12538
rect 3032 12486 3044 12538
rect 3044 12486 3058 12538
rect 3082 12486 3096 12538
rect 3096 12486 3108 12538
rect 3108 12486 3138 12538
rect 3162 12486 3172 12538
rect 3172 12486 3218 12538
rect 2922 12484 2978 12486
rect 3002 12484 3058 12486
rect 3082 12484 3138 12486
rect 3162 12484 3218 12486
rect 2922 11450 2978 11452
rect 3002 11450 3058 11452
rect 3082 11450 3138 11452
rect 3162 11450 3218 11452
rect 2922 11398 2968 11450
rect 2968 11398 2978 11450
rect 3002 11398 3032 11450
rect 3032 11398 3044 11450
rect 3044 11398 3058 11450
rect 3082 11398 3096 11450
rect 3096 11398 3108 11450
rect 3108 11398 3138 11450
rect 3162 11398 3172 11450
rect 3172 11398 3218 11450
rect 2922 11396 2978 11398
rect 3002 11396 3058 11398
rect 3082 11396 3138 11398
rect 3162 11396 3218 11398
rect 4888 15258 4944 15260
rect 4968 15258 5024 15260
rect 5048 15258 5104 15260
rect 5128 15258 5184 15260
rect 4888 15206 4934 15258
rect 4934 15206 4944 15258
rect 4968 15206 4998 15258
rect 4998 15206 5010 15258
rect 5010 15206 5024 15258
rect 5048 15206 5062 15258
rect 5062 15206 5074 15258
rect 5074 15206 5104 15258
rect 5128 15206 5138 15258
rect 5138 15206 5184 15258
rect 4888 15204 4944 15206
rect 4968 15204 5024 15206
rect 5048 15204 5104 15206
rect 5128 15204 5184 15206
rect 5722 15000 5778 15056
rect 4888 14170 4944 14172
rect 4968 14170 5024 14172
rect 5048 14170 5104 14172
rect 5128 14170 5184 14172
rect 4888 14118 4934 14170
rect 4934 14118 4944 14170
rect 4968 14118 4998 14170
rect 4998 14118 5010 14170
rect 5010 14118 5024 14170
rect 5048 14118 5062 14170
rect 5062 14118 5074 14170
rect 5074 14118 5104 14170
rect 5128 14118 5138 14170
rect 5138 14118 5184 14170
rect 4888 14116 4944 14118
rect 4968 14116 5024 14118
rect 5048 14116 5104 14118
rect 5128 14116 5184 14118
rect 4066 13912 4122 13968
rect 2922 10362 2978 10364
rect 3002 10362 3058 10364
rect 3082 10362 3138 10364
rect 3162 10362 3218 10364
rect 2922 10310 2968 10362
rect 2968 10310 2978 10362
rect 3002 10310 3032 10362
rect 3032 10310 3044 10362
rect 3044 10310 3058 10362
rect 3082 10310 3096 10362
rect 3096 10310 3108 10362
rect 3108 10310 3138 10362
rect 3162 10310 3172 10362
rect 3172 10310 3218 10362
rect 2922 10308 2978 10310
rect 3002 10308 3058 10310
rect 3082 10308 3138 10310
rect 3162 10308 3218 10310
rect 5630 13932 5686 13968
rect 5630 13912 5632 13932
rect 5632 13912 5684 13932
rect 5684 13912 5686 13932
rect 4888 13082 4944 13084
rect 4968 13082 5024 13084
rect 5048 13082 5104 13084
rect 5128 13082 5184 13084
rect 4888 13030 4934 13082
rect 4934 13030 4944 13082
rect 4968 13030 4998 13082
rect 4998 13030 5010 13082
rect 5010 13030 5024 13082
rect 5048 13030 5062 13082
rect 5062 13030 5074 13082
rect 5074 13030 5104 13082
rect 5128 13030 5138 13082
rect 5138 13030 5184 13082
rect 4888 13028 4944 13030
rect 4968 13028 5024 13030
rect 5048 13028 5104 13030
rect 5128 13028 5184 13030
rect 2922 9274 2978 9276
rect 3002 9274 3058 9276
rect 3082 9274 3138 9276
rect 3162 9274 3218 9276
rect 2922 9222 2968 9274
rect 2968 9222 2978 9274
rect 3002 9222 3032 9274
rect 3032 9222 3044 9274
rect 3044 9222 3058 9274
rect 3082 9222 3096 9274
rect 3096 9222 3108 9274
rect 3108 9222 3138 9274
rect 3162 9222 3172 9274
rect 3172 9222 3218 9274
rect 2922 9220 2978 9222
rect 3002 9220 3058 9222
rect 3082 9220 3138 9222
rect 3162 9220 3218 9222
rect 2922 8186 2978 8188
rect 3002 8186 3058 8188
rect 3082 8186 3138 8188
rect 3162 8186 3218 8188
rect 2922 8134 2968 8186
rect 2968 8134 2978 8186
rect 3002 8134 3032 8186
rect 3032 8134 3044 8186
rect 3044 8134 3058 8186
rect 3082 8134 3096 8186
rect 3096 8134 3108 8186
rect 3108 8134 3138 8186
rect 3162 8134 3172 8186
rect 3172 8134 3218 8186
rect 2922 8132 2978 8134
rect 3002 8132 3058 8134
rect 3082 8132 3138 8134
rect 3162 8132 3218 8134
rect 2922 7098 2978 7100
rect 3002 7098 3058 7100
rect 3082 7098 3138 7100
rect 3162 7098 3218 7100
rect 2922 7046 2968 7098
rect 2968 7046 2978 7098
rect 3002 7046 3032 7098
rect 3032 7046 3044 7098
rect 3044 7046 3058 7098
rect 3082 7046 3096 7098
rect 3096 7046 3108 7098
rect 3108 7046 3138 7098
rect 3162 7046 3172 7098
rect 3172 7046 3218 7098
rect 2922 7044 2978 7046
rect 3002 7044 3058 7046
rect 3082 7044 3138 7046
rect 3162 7044 3218 7046
rect 4888 11994 4944 11996
rect 4968 11994 5024 11996
rect 5048 11994 5104 11996
rect 5128 11994 5184 11996
rect 4888 11942 4934 11994
rect 4934 11942 4944 11994
rect 4968 11942 4998 11994
rect 4998 11942 5010 11994
rect 5010 11942 5024 11994
rect 5048 11942 5062 11994
rect 5062 11942 5074 11994
rect 5074 11942 5104 11994
rect 5128 11942 5138 11994
rect 5138 11942 5184 11994
rect 4888 11940 4944 11942
rect 4968 11940 5024 11942
rect 5048 11940 5104 11942
rect 5128 11940 5184 11942
rect 4888 10906 4944 10908
rect 4968 10906 5024 10908
rect 5048 10906 5104 10908
rect 5128 10906 5184 10908
rect 4888 10854 4934 10906
rect 4934 10854 4944 10906
rect 4968 10854 4998 10906
rect 4998 10854 5010 10906
rect 5010 10854 5024 10906
rect 5048 10854 5062 10906
rect 5062 10854 5074 10906
rect 5074 10854 5104 10906
rect 5128 10854 5138 10906
rect 5138 10854 5184 10906
rect 4888 10852 4944 10854
rect 4968 10852 5024 10854
rect 5048 10852 5104 10854
rect 5128 10852 5184 10854
rect 6550 15020 6606 15056
rect 6550 15000 6552 15020
rect 6552 15000 6604 15020
rect 6604 15000 6606 15020
rect 6855 14714 6911 14716
rect 6935 14714 6991 14716
rect 7015 14714 7071 14716
rect 7095 14714 7151 14716
rect 6855 14662 6901 14714
rect 6901 14662 6911 14714
rect 6935 14662 6965 14714
rect 6965 14662 6977 14714
rect 6977 14662 6991 14714
rect 7015 14662 7029 14714
rect 7029 14662 7041 14714
rect 7041 14662 7071 14714
rect 7095 14662 7105 14714
rect 7105 14662 7151 14714
rect 6855 14660 6911 14662
rect 6935 14660 6991 14662
rect 7015 14660 7071 14662
rect 7095 14660 7151 14662
rect 8821 15258 8877 15260
rect 8901 15258 8957 15260
rect 8981 15258 9037 15260
rect 9061 15258 9117 15260
rect 8821 15206 8867 15258
rect 8867 15206 8877 15258
rect 8901 15206 8931 15258
rect 8931 15206 8943 15258
rect 8943 15206 8957 15258
rect 8981 15206 8995 15258
rect 8995 15206 9007 15258
rect 9007 15206 9037 15258
rect 9061 15206 9071 15258
rect 9071 15206 9117 15258
rect 8821 15204 8877 15206
rect 8901 15204 8957 15206
rect 8981 15204 9037 15206
rect 9061 15204 9117 15206
rect 12754 15258 12810 15260
rect 12834 15258 12890 15260
rect 12914 15258 12970 15260
rect 12994 15258 13050 15260
rect 12754 15206 12800 15258
rect 12800 15206 12810 15258
rect 12834 15206 12864 15258
rect 12864 15206 12876 15258
rect 12876 15206 12890 15258
rect 12914 15206 12928 15258
rect 12928 15206 12940 15258
rect 12940 15206 12970 15258
rect 12994 15206 13004 15258
rect 13004 15206 13050 15258
rect 12754 15204 12810 15206
rect 12834 15204 12890 15206
rect 12914 15204 12970 15206
rect 12994 15204 13050 15206
rect 10788 14714 10844 14716
rect 10868 14714 10924 14716
rect 10948 14714 11004 14716
rect 11028 14714 11084 14716
rect 10788 14662 10834 14714
rect 10834 14662 10844 14714
rect 10868 14662 10898 14714
rect 10898 14662 10910 14714
rect 10910 14662 10924 14714
rect 10948 14662 10962 14714
rect 10962 14662 10974 14714
rect 10974 14662 11004 14714
rect 11028 14662 11038 14714
rect 11038 14662 11084 14714
rect 10788 14660 10844 14662
rect 10868 14660 10924 14662
rect 10948 14660 11004 14662
rect 11028 14660 11084 14662
rect 6855 13626 6911 13628
rect 6935 13626 6991 13628
rect 7015 13626 7071 13628
rect 7095 13626 7151 13628
rect 6855 13574 6901 13626
rect 6901 13574 6911 13626
rect 6935 13574 6965 13626
rect 6965 13574 6977 13626
rect 6977 13574 6991 13626
rect 7015 13574 7029 13626
rect 7029 13574 7041 13626
rect 7041 13574 7071 13626
rect 7095 13574 7105 13626
rect 7105 13574 7151 13626
rect 6855 13572 6911 13574
rect 6935 13572 6991 13574
rect 7015 13572 7071 13574
rect 7095 13572 7151 13574
rect 8821 14170 8877 14172
rect 8901 14170 8957 14172
rect 8981 14170 9037 14172
rect 9061 14170 9117 14172
rect 8821 14118 8867 14170
rect 8867 14118 8877 14170
rect 8901 14118 8931 14170
rect 8931 14118 8943 14170
rect 8943 14118 8957 14170
rect 8981 14118 8995 14170
rect 8995 14118 9007 14170
rect 9007 14118 9037 14170
rect 9061 14118 9071 14170
rect 9071 14118 9117 14170
rect 8821 14116 8877 14118
rect 8901 14116 8957 14118
rect 8981 14116 9037 14118
rect 9061 14116 9117 14118
rect 12754 14170 12810 14172
rect 12834 14170 12890 14172
rect 12914 14170 12970 14172
rect 12994 14170 13050 14172
rect 12754 14118 12800 14170
rect 12800 14118 12810 14170
rect 12834 14118 12864 14170
rect 12864 14118 12876 14170
rect 12876 14118 12890 14170
rect 12914 14118 12928 14170
rect 12928 14118 12940 14170
rect 12940 14118 12970 14170
rect 12994 14118 13004 14170
rect 13004 14118 13050 14170
rect 12754 14116 12810 14118
rect 12834 14116 12890 14118
rect 12914 14116 12970 14118
rect 12994 14116 13050 14118
rect 7838 13912 7894 13968
rect 10788 13626 10844 13628
rect 10868 13626 10924 13628
rect 10948 13626 11004 13628
rect 11028 13626 11084 13628
rect 10788 13574 10834 13626
rect 10834 13574 10844 13626
rect 10868 13574 10898 13626
rect 10898 13574 10910 13626
rect 10910 13574 10924 13626
rect 10948 13574 10962 13626
rect 10962 13574 10974 13626
rect 10974 13574 11004 13626
rect 11028 13574 11038 13626
rect 11038 13574 11084 13626
rect 10788 13572 10844 13574
rect 10868 13572 10924 13574
rect 10948 13572 11004 13574
rect 11028 13572 11084 13574
rect 8821 13082 8877 13084
rect 8901 13082 8957 13084
rect 8981 13082 9037 13084
rect 9061 13082 9117 13084
rect 8821 13030 8867 13082
rect 8867 13030 8877 13082
rect 8901 13030 8931 13082
rect 8931 13030 8943 13082
rect 8943 13030 8957 13082
rect 8981 13030 8995 13082
rect 8995 13030 9007 13082
rect 9007 13030 9037 13082
rect 9061 13030 9071 13082
rect 9071 13030 9117 13082
rect 8821 13028 8877 13030
rect 8901 13028 8957 13030
rect 8981 13028 9037 13030
rect 9061 13028 9117 13030
rect 12754 13082 12810 13084
rect 12834 13082 12890 13084
rect 12914 13082 12970 13084
rect 12994 13082 13050 13084
rect 12754 13030 12800 13082
rect 12800 13030 12810 13082
rect 12834 13030 12864 13082
rect 12864 13030 12876 13082
rect 12876 13030 12890 13082
rect 12914 13030 12928 13082
rect 12928 13030 12940 13082
rect 12940 13030 12970 13082
rect 12994 13030 13004 13082
rect 13004 13030 13050 13082
rect 12754 13028 12810 13030
rect 12834 13028 12890 13030
rect 12914 13028 12970 13030
rect 12994 13028 13050 13030
rect 6855 12538 6911 12540
rect 6935 12538 6991 12540
rect 7015 12538 7071 12540
rect 7095 12538 7151 12540
rect 6855 12486 6901 12538
rect 6901 12486 6911 12538
rect 6935 12486 6965 12538
rect 6965 12486 6977 12538
rect 6977 12486 6991 12538
rect 7015 12486 7029 12538
rect 7029 12486 7041 12538
rect 7041 12486 7071 12538
rect 7095 12486 7105 12538
rect 7105 12486 7151 12538
rect 6855 12484 6911 12486
rect 6935 12484 6991 12486
rect 7015 12484 7071 12486
rect 7095 12484 7151 12486
rect 6855 11450 6911 11452
rect 6935 11450 6991 11452
rect 7015 11450 7071 11452
rect 7095 11450 7151 11452
rect 6855 11398 6901 11450
rect 6901 11398 6911 11450
rect 6935 11398 6965 11450
rect 6965 11398 6977 11450
rect 6977 11398 6991 11450
rect 7015 11398 7029 11450
rect 7029 11398 7041 11450
rect 7041 11398 7071 11450
rect 7095 11398 7105 11450
rect 7105 11398 7151 11450
rect 6855 11396 6911 11398
rect 6935 11396 6991 11398
rect 7015 11396 7071 11398
rect 7095 11396 7151 11398
rect 6855 10362 6911 10364
rect 6935 10362 6991 10364
rect 7015 10362 7071 10364
rect 7095 10362 7151 10364
rect 6855 10310 6901 10362
rect 6901 10310 6911 10362
rect 6935 10310 6965 10362
rect 6965 10310 6977 10362
rect 6977 10310 6991 10362
rect 7015 10310 7029 10362
rect 7029 10310 7041 10362
rect 7041 10310 7071 10362
rect 7095 10310 7105 10362
rect 7105 10310 7151 10362
rect 6855 10308 6911 10310
rect 6935 10308 6991 10310
rect 7015 10308 7071 10310
rect 7095 10308 7151 10310
rect 10788 12538 10844 12540
rect 10868 12538 10924 12540
rect 10948 12538 11004 12540
rect 11028 12538 11084 12540
rect 10788 12486 10834 12538
rect 10834 12486 10844 12538
rect 10868 12486 10898 12538
rect 10898 12486 10910 12538
rect 10910 12486 10924 12538
rect 10948 12486 10962 12538
rect 10962 12486 10974 12538
rect 10974 12486 11004 12538
rect 11028 12486 11038 12538
rect 11038 12486 11084 12538
rect 10788 12484 10844 12486
rect 10868 12484 10924 12486
rect 10948 12484 11004 12486
rect 11028 12484 11084 12486
rect 8821 11994 8877 11996
rect 8901 11994 8957 11996
rect 8981 11994 9037 11996
rect 9061 11994 9117 11996
rect 8821 11942 8867 11994
rect 8867 11942 8877 11994
rect 8901 11942 8931 11994
rect 8931 11942 8943 11994
rect 8943 11942 8957 11994
rect 8981 11942 8995 11994
rect 8995 11942 9007 11994
rect 9007 11942 9037 11994
rect 9061 11942 9071 11994
rect 9071 11942 9117 11994
rect 8821 11940 8877 11942
rect 8901 11940 8957 11942
rect 8981 11940 9037 11942
rect 9061 11940 9117 11942
rect 12754 11994 12810 11996
rect 12834 11994 12890 11996
rect 12914 11994 12970 11996
rect 12994 11994 13050 11996
rect 12754 11942 12800 11994
rect 12800 11942 12810 11994
rect 12834 11942 12864 11994
rect 12864 11942 12876 11994
rect 12876 11942 12890 11994
rect 12914 11942 12928 11994
rect 12928 11942 12940 11994
rect 12940 11942 12970 11994
rect 12994 11942 13004 11994
rect 13004 11942 13050 11994
rect 12754 11940 12810 11942
rect 12834 11940 12890 11942
rect 12914 11940 12970 11942
rect 12994 11940 13050 11942
rect 8821 10906 8877 10908
rect 8901 10906 8957 10908
rect 8981 10906 9037 10908
rect 9061 10906 9117 10908
rect 8821 10854 8867 10906
rect 8867 10854 8877 10906
rect 8901 10854 8931 10906
rect 8931 10854 8943 10906
rect 8943 10854 8957 10906
rect 8981 10854 8995 10906
rect 8995 10854 9007 10906
rect 9007 10854 9037 10906
rect 9061 10854 9071 10906
rect 9071 10854 9117 10906
rect 8821 10852 8877 10854
rect 8901 10852 8957 10854
rect 8981 10852 9037 10854
rect 9061 10852 9117 10854
rect 10788 11450 10844 11452
rect 10868 11450 10924 11452
rect 10948 11450 11004 11452
rect 11028 11450 11084 11452
rect 10788 11398 10834 11450
rect 10834 11398 10844 11450
rect 10868 11398 10898 11450
rect 10898 11398 10910 11450
rect 10910 11398 10924 11450
rect 10948 11398 10962 11450
rect 10962 11398 10974 11450
rect 10974 11398 11004 11450
rect 11028 11398 11038 11450
rect 11038 11398 11084 11450
rect 10788 11396 10844 11398
rect 10868 11396 10924 11398
rect 10948 11396 11004 11398
rect 11028 11396 11084 11398
rect 14721 15802 14777 15804
rect 14801 15802 14857 15804
rect 14881 15802 14937 15804
rect 14961 15802 15017 15804
rect 14721 15750 14767 15802
rect 14767 15750 14777 15802
rect 14801 15750 14831 15802
rect 14831 15750 14843 15802
rect 14843 15750 14857 15802
rect 14881 15750 14895 15802
rect 14895 15750 14907 15802
rect 14907 15750 14937 15802
rect 14961 15750 14971 15802
rect 14971 15750 15017 15802
rect 14721 15748 14777 15750
rect 14801 15748 14857 15750
rect 14881 15748 14937 15750
rect 14961 15748 15017 15750
rect 16687 15258 16743 15260
rect 16767 15258 16823 15260
rect 16847 15258 16903 15260
rect 16927 15258 16983 15260
rect 16687 15206 16733 15258
rect 16733 15206 16743 15258
rect 16767 15206 16797 15258
rect 16797 15206 16809 15258
rect 16809 15206 16823 15258
rect 16847 15206 16861 15258
rect 16861 15206 16873 15258
rect 16873 15206 16903 15258
rect 16927 15206 16937 15258
rect 16937 15206 16983 15258
rect 16687 15204 16743 15206
rect 16767 15204 16823 15206
rect 16847 15204 16903 15206
rect 16927 15204 16983 15206
rect 14721 14714 14777 14716
rect 14801 14714 14857 14716
rect 14881 14714 14937 14716
rect 14961 14714 15017 14716
rect 14721 14662 14767 14714
rect 14767 14662 14777 14714
rect 14801 14662 14831 14714
rect 14831 14662 14843 14714
rect 14843 14662 14857 14714
rect 14881 14662 14895 14714
rect 14895 14662 14907 14714
rect 14907 14662 14937 14714
rect 14961 14662 14971 14714
rect 14971 14662 15017 14714
rect 14721 14660 14777 14662
rect 14801 14660 14857 14662
rect 14881 14660 14937 14662
rect 14961 14660 15017 14662
rect 16687 14170 16743 14172
rect 16767 14170 16823 14172
rect 16847 14170 16903 14172
rect 16927 14170 16983 14172
rect 16687 14118 16733 14170
rect 16733 14118 16743 14170
rect 16767 14118 16797 14170
rect 16797 14118 16809 14170
rect 16809 14118 16823 14170
rect 16847 14118 16861 14170
rect 16861 14118 16873 14170
rect 16873 14118 16903 14170
rect 16927 14118 16937 14170
rect 16937 14118 16983 14170
rect 16687 14116 16743 14118
rect 16767 14116 16823 14118
rect 16847 14116 16903 14118
rect 16927 14116 16983 14118
rect 14721 13626 14777 13628
rect 14801 13626 14857 13628
rect 14881 13626 14937 13628
rect 14961 13626 15017 13628
rect 14721 13574 14767 13626
rect 14767 13574 14777 13626
rect 14801 13574 14831 13626
rect 14831 13574 14843 13626
rect 14843 13574 14857 13626
rect 14881 13574 14895 13626
rect 14895 13574 14907 13626
rect 14907 13574 14937 13626
rect 14961 13574 14971 13626
rect 14971 13574 15017 13626
rect 14721 13572 14777 13574
rect 14801 13572 14857 13574
rect 14881 13572 14937 13574
rect 14961 13572 15017 13574
rect 16687 13082 16743 13084
rect 16767 13082 16823 13084
rect 16847 13082 16903 13084
rect 16927 13082 16983 13084
rect 16687 13030 16733 13082
rect 16733 13030 16743 13082
rect 16767 13030 16797 13082
rect 16797 13030 16809 13082
rect 16809 13030 16823 13082
rect 16847 13030 16861 13082
rect 16861 13030 16873 13082
rect 16873 13030 16903 13082
rect 16927 13030 16937 13082
rect 16937 13030 16983 13082
rect 16687 13028 16743 13030
rect 16767 13028 16823 13030
rect 16847 13028 16903 13030
rect 16927 13028 16983 13030
rect 14721 12538 14777 12540
rect 14801 12538 14857 12540
rect 14881 12538 14937 12540
rect 14961 12538 15017 12540
rect 14721 12486 14767 12538
rect 14767 12486 14777 12538
rect 14801 12486 14831 12538
rect 14831 12486 14843 12538
rect 14843 12486 14857 12538
rect 14881 12486 14895 12538
rect 14895 12486 14907 12538
rect 14907 12486 14937 12538
rect 14961 12486 14971 12538
rect 14971 12486 15017 12538
rect 14721 12484 14777 12486
rect 14801 12484 14857 12486
rect 14881 12484 14937 12486
rect 14961 12484 15017 12486
rect 16687 11994 16743 11996
rect 16767 11994 16823 11996
rect 16847 11994 16903 11996
rect 16927 11994 16983 11996
rect 16687 11942 16733 11994
rect 16733 11942 16743 11994
rect 16767 11942 16797 11994
rect 16797 11942 16809 11994
rect 16809 11942 16823 11994
rect 16847 11942 16861 11994
rect 16861 11942 16873 11994
rect 16873 11942 16903 11994
rect 16927 11942 16937 11994
rect 16937 11942 16983 11994
rect 16687 11940 16743 11942
rect 16767 11940 16823 11942
rect 16847 11940 16903 11942
rect 16927 11940 16983 11942
rect 14721 11450 14777 11452
rect 14801 11450 14857 11452
rect 14881 11450 14937 11452
rect 14961 11450 15017 11452
rect 14721 11398 14767 11450
rect 14767 11398 14777 11450
rect 14801 11398 14831 11450
rect 14831 11398 14843 11450
rect 14843 11398 14857 11450
rect 14881 11398 14895 11450
rect 14895 11398 14907 11450
rect 14907 11398 14937 11450
rect 14961 11398 14971 11450
rect 14971 11398 15017 11450
rect 14721 11396 14777 11398
rect 14801 11396 14857 11398
rect 14881 11396 14937 11398
rect 14961 11396 15017 11398
rect 12754 10906 12810 10908
rect 12834 10906 12890 10908
rect 12914 10906 12970 10908
rect 12994 10906 13050 10908
rect 12754 10854 12800 10906
rect 12800 10854 12810 10906
rect 12834 10854 12864 10906
rect 12864 10854 12876 10906
rect 12876 10854 12890 10906
rect 12914 10854 12928 10906
rect 12928 10854 12940 10906
rect 12940 10854 12970 10906
rect 12994 10854 13004 10906
rect 13004 10854 13050 10906
rect 12754 10852 12810 10854
rect 12834 10852 12890 10854
rect 12914 10852 12970 10854
rect 12994 10852 13050 10854
rect 16687 10906 16743 10908
rect 16767 10906 16823 10908
rect 16847 10906 16903 10908
rect 16927 10906 16983 10908
rect 16687 10854 16733 10906
rect 16733 10854 16743 10906
rect 16767 10854 16797 10906
rect 16797 10854 16809 10906
rect 16809 10854 16823 10906
rect 16847 10854 16861 10906
rect 16861 10854 16873 10906
rect 16873 10854 16903 10906
rect 16927 10854 16937 10906
rect 16937 10854 16983 10906
rect 16687 10852 16743 10854
rect 16767 10852 16823 10854
rect 16847 10852 16903 10854
rect 16927 10852 16983 10854
rect 10788 10362 10844 10364
rect 10868 10362 10924 10364
rect 10948 10362 11004 10364
rect 11028 10362 11084 10364
rect 10788 10310 10834 10362
rect 10834 10310 10844 10362
rect 10868 10310 10898 10362
rect 10898 10310 10910 10362
rect 10910 10310 10924 10362
rect 10948 10310 10962 10362
rect 10962 10310 10974 10362
rect 10974 10310 11004 10362
rect 11028 10310 11038 10362
rect 11038 10310 11084 10362
rect 10788 10308 10844 10310
rect 10868 10308 10924 10310
rect 10948 10308 11004 10310
rect 11028 10308 11084 10310
rect 14721 10362 14777 10364
rect 14801 10362 14857 10364
rect 14881 10362 14937 10364
rect 14961 10362 15017 10364
rect 14721 10310 14767 10362
rect 14767 10310 14777 10362
rect 14801 10310 14831 10362
rect 14831 10310 14843 10362
rect 14843 10310 14857 10362
rect 14881 10310 14895 10362
rect 14895 10310 14907 10362
rect 14907 10310 14937 10362
rect 14961 10310 14971 10362
rect 14971 10310 15017 10362
rect 14721 10308 14777 10310
rect 14801 10308 14857 10310
rect 14881 10308 14937 10310
rect 14961 10308 15017 10310
rect 4888 9818 4944 9820
rect 4968 9818 5024 9820
rect 5048 9818 5104 9820
rect 5128 9818 5184 9820
rect 4888 9766 4934 9818
rect 4934 9766 4944 9818
rect 4968 9766 4998 9818
rect 4998 9766 5010 9818
rect 5010 9766 5024 9818
rect 5048 9766 5062 9818
rect 5062 9766 5074 9818
rect 5074 9766 5104 9818
rect 5128 9766 5138 9818
rect 5138 9766 5184 9818
rect 4888 9764 4944 9766
rect 4968 9764 5024 9766
rect 5048 9764 5104 9766
rect 5128 9764 5184 9766
rect 8821 9818 8877 9820
rect 8901 9818 8957 9820
rect 8981 9818 9037 9820
rect 9061 9818 9117 9820
rect 8821 9766 8867 9818
rect 8867 9766 8877 9818
rect 8901 9766 8931 9818
rect 8931 9766 8943 9818
rect 8943 9766 8957 9818
rect 8981 9766 8995 9818
rect 8995 9766 9007 9818
rect 9007 9766 9037 9818
rect 9061 9766 9071 9818
rect 9071 9766 9117 9818
rect 8821 9764 8877 9766
rect 8901 9764 8957 9766
rect 8981 9764 9037 9766
rect 9061 9764 9117 9766
rect 12754 9818 12810 9820
rect 12834 9818 12890 9820
rect 12914 9818 12970 9820
rect 12994 9818 13050 9820
rect 12754 9766 12800 9818
rect 12800 9766 12810 9818
rect 12834 9766 12864 9818
rect 12864 9766 12876 9818
rect 12876 9766 12890 9818
rect 12914 9766 12928 9818
rect 12928 9766 12940 9818
rect 12940 9766 12970 9818
rect 12994 9766 13004 9818
rect 13004 9766 13050 9818
rect 12754 9764 12810 9766
rect 12834 9764 12890 9766
rect 12914 9764 12970 9766
rect 12994 9764 13050 9766
rect 16687 9818 16743 9820
rect 16767 9818 16823 9820
rect 16847 9818 16903 9820
rect 16927 9818 16983 9820
rect 16687 9766 16733 9818
rect 16733 9766 16743 9818
rect 16767 9766 16797 9818
rect 16797 9766 16809 9818
rect 16809 9766 16823 9818
rect 16847 9766 16861 9818
rect 16861 9766 16873 9818
rect 16873 9766 16903 9818
rect 16927 9766 16937 9818
rect 16937 9766 16983 9818
rect 16687 9764 16743 9766
rect 16767 9764 16823 9766
rect 16847 9764 16903 9766
rect 16927 9764 16983 9766
rect 6855 9274 6911 9276
rect 6935 9274 6991 9276
rect 7015 9274 7071 9276
rect 7095 9274 7151 9276
rect 6855 9222 6901 9274
rect 6901 9222 6911 9274
rect 6935 9222 6965 9274
rect 6965 9222 6977 9274
rect 6977 9222 6991 9274
rect 7015 9222 7029 9274
rect 7029 9222 7041 9274
rect 7041 9222 7071 9274
rect 7095 9222 7105 9274
rect 7105 9222 7151 9274
rect 6855 9220 6911 9222
rect 6935 9220 6991 9222
rect 7015 9220 7071 9222
rect 7095 9220 7151 9222
rect 10788 9274 10844 9276
rect 10868 9274 10924 9276
rect 10948 9274 11004 9276
rect 11028 9274 11084 9276
rect 10788 9222 10834 9274
rect 10834 9222 10844 9274
rect 10868 9222 10898 9274
rect 10898 9222 10910 9274
rect 10910 9222 10924 9274
rect 10948 9222 10962 9274
rect 10962 9222 10974 9274
rect 10974 9222 11004 9274
rect 11028 9222 11038 9274
rect 11038 9222 11084 9274
rect 10788 9220 10844 9222
rect 10868 9220 10924 9222
rect 10948 9220 11004 9222
rect 11028 9220 11084 9222
rect 14721 9274 14777 9276
rect 14801 9274 14857 9276
rect 14881 9274 14937 9276
rect 14961 9274 15017 9276
rect 14721 9222 14767 9274
rect 14767 9222 14777 9274
rect 14801 9222 14831 9274
rect 14831 9222 14843 9274
rect 14843 9222 14857 9274
rect 14881 9222 14895 9274
rect 14895 9222 14907 9274
rect 14907 9222 14937 9274
rect 14961 9222 14971 9274
rect 14971 9222 15017 9274
rect 14721 9220 14777 9222
rect 14801 9220 14857 9222
rect 14881 9220 14937 9222
rect 14961 9220 15017 9222
rect 4888 8730 4944 8732
rect 4968 8730 5024 8732
rect 5048 8730 5104 8732
rect 5128 8730 5184 8732
rect 4888 8678 4934 8730
rect 4934 8678 4944 8730
rect 4968 8678 4998 8730
rect 4998 8678 5010 8730
rect 5010 8678 5024 8730
rect 5048 8678 5062 8730
rect 5062 8678 5074 8730
rect 5074 8678 5104 8730
rect 5128 8678 5138 8730
rect 5138 8678 5184 8730
rect 4888 8676 4944 8678
rect 4968 8676 5024 8678
rect 5048 8676 5104 8678
rect 5128 8676 5184 8678
rect 8821 8730 8877 8732
rect 8901 8730 8957 8732
rect 8981 8730 9037 8732
rect 9061 8730 9117 8732
rect 8821 8678 8867 8730
rect 8867 8678 8877 8730
rect 8901 8678 8931 8730
rect 8931 8678 8943 8730
rect 8943 8678 8957 8730
rect 8981 8678 8995 8730
rect 8995 8678 9007 8730
rect 9007 8678 9037 8730
rect 9061 8678 9071 8730
rect 9071 8678 9117 8730
rect 8821 8676 8877 8678
rect 8901 8676 8957 8678
rect 8981 8676 9037 8678
rect 9061 8676 9117 8678
rect 12754 8730 12810 8732
rect 12834 8730 12890 8732
rect 12914 8730 12970 8732
rect 12994 8730 13050 8732
rect 12754 8678 12800 8730
rect 12800 8678 12810 8730
rect 12834 8678 12864 8730
rect 12864 8678 12876 8730
rect 12876 8678 12890 8730
rect 12914 8678 12928 8730
rect 12928 8678 12940 8730
rect 12940 8678 12970 8730
rect 12994 8678 13004 8730
rect 13004 8678 13050 8730
rect 12754 8676 12810 8678
rect 12834 8676 12890 8678
rect 12914 8676 12970 8678
rect 12994 8676 13050 8678
rect 16687 8730 16743 8732
rect 16767 8730 16823 8732
rect 16847 8730 16903 8732
rect 16927 8730 16983 8732
rect 16687 8678 16733 8730
rect 16733 8678 16743 8730
rect 16767 8678 16797 8730
rect 16797 8678 16809 8730
rect 16809 8678 16823 8730
rect 16847 8678 16861 8730
rect 16861 8678 16873 8730
rect 16873 8678 16903 8730
rect 16927 8678 16937 8730
rect 16937 8678 16983 8730
rect 16687 8676 16743 8678
rect 16767 8676 16823 8678
rect 16847 8676 16903 8678
rect 16927 8676 16983 8678
rect 6855 8186 6911 8188
rect 6935 8186 6991 8188
rect 7015 8186 7071 8188
rect 7095 8186 7151 8188
rect 6855 8134 6901 8186
rect 6901 8134 6911 8186
rect 6935 8134 6965 8186
rect 6965 8134 6977 8186
rect 6977 8134 6991 8186
rect 7015 8134 7029 8186
rect 7029 8134 7041 8186
rect 7041 8134 7071 8186
rect 7095 8134 7105 8186
rect 7105 8134 7151 8186
rect 6855 8132 6911 8134
rect 6935 8132 6991 8134
rect 7015 8132 7071 8134
rect 7095 8132 7151 8134
rect 10788 8186 10844 8188
rect 10868 8186 10924 8188
rect 10948 8186 11004 8188
rect 11028 8186 11084 8188
rect 10788 8134 10834 8186
rect 10834 8134 10844 8186
rect 10868 8134 10898 8186
rect 10898 8134 10910 8186
rect 10910 8134 10924 8186
rect 10948 8134 10962 8186
rect 10962 8134 10974 8186
rect 10974 8134 11004 8186
rect 11028 8134 11038 8186
rect 11038 8134 11084 8186
rect 10788 8132 10844 8134
rect 10868 8132 10924 8134
rect 10948 8132 11004 8134
rect 11028 8132 11084 8134
rect 14721 8186 14777 8188
rect 14801 8186 14857 8188
rect 14881 8186 14937 8188
rect 14961 8186 15017 8188
rect 14721 8134 14767 8186
rect 14767 8134 14777 8186
rect 14801 8134 14831 8186
rect 14831 8134 14843 8186
rect 14843 8134 14857 8186
rect 14881 8134 14895 8186
rect 14895 8134 14907 8186
rect 14907 8134 14937 8186
rect 14961 8134 14971 8186
rect 14971 8134 15017 8186
rect 14721 8132 14777 8134
rect 14801 8132 14857 8134
rect 14881 8132 14937 8134
rect 14961 8132 15017 8134
rect 4888 7642 4944 7644
rect 4968 7642 5024 7644
rect 5048 7642 5104 7644
rect 5128 7642 5184 7644
rect 4888 7590 4934 7642
rect 4934 7590 4944 7642
rect 4968 7590 4998 7642
rect 4998 7590 5010 7642
rect 5010 7590 5024 7642
rect 5048 7590 5062 7642
rect 5062 7590 5074 7642
rect 5074 7590 5104 7642
rect 5128 7590 5138 7642
rect 5138 7590 5184 7642
rect 4888 7588 4944 7590
rect 4968 7588 5024 7590
rect 5048 7588 5104 7590
rect 5128 7588 5184 7590
rect 8821 7642 8877 7644
rect 8901 7642 8957 7644
rect 8981 7642 9037 7644
rect 9061 7642 9117 7644
rect 8821 7590 8867 7642
rect 8867 7590 8877 7642
rect 8901 7590 8931 7642
rect 8931 7590 8943 7642
rect 8943 7590 8957 7642
rect 8981 7590 8995 7642
rect 8995 7590 9007 7642
rect 9007 7590 9037 7642
rect 9061 7590 9071 7642
rect 9071 7590 9117 7642
rect 8821 7588 8877 7590
rect 8901 7588 8957 7590
rect 8981 7588 9037 7590
rect 9061 7588 9117 7590
rect 12754 7642 12810 7644
rect 12834 7642 12890 7644
rect 12914 7642 12970 7644
rect 12994 7642 13050 7644
rect 12754 7590 12800 7642
rect 12800 7590 12810 7642
rect 12834 7590 12864 7642
rect 12864 7590 12876 7642
rect 12876 7590 12890 7642
rect 12914 7590 12928 7642
rect 12928 7590 12940 7642
rect 12940 7590 12970 7642
rect 12994 7590 13004 7642
rect 13004 7590 13050 7642
rect 12754 7588 12810 7590
rect 12834 7588 12890 7590
rect 12914 7588 12970 7590
rect 12994 7588 13050 7590
rect 16687 7642 16743 7644
rect 16767 7642 16823 7644
rect 16847 7642 16903 7644
rect 16927 7642 16983 7644
rect 16687 7590 16733 7642
rect 16733 7590 16743 7642
rect 16767 7590 16797 7642
rect 16797 7590 16809 7642
rect 16809 7590 16823 7642
rect 16847 7590 16861 7642
rect 16861 7590 16873 7642
rect 16873 7590 16903 7642
rect 16927 7590 16937 7642
rect 16937 7590 16983 7642
rect 16687 7588 16743 7590
rect 16767 7588 16823 7590
rect 16847 7588 16903 7590
rect 16927 7588 16983 7590
rect 6855 7098 6911 7100
rect 6935 7098 6991 7100
rect 7015 7098 7071 7100
rect 7095 7098 7151 7100
rect 6855 7046 6901 7098
rect 6901 7046 6911 7098
rect 6935 7046 6965 7098
rect 6965 7046 6977 7098
rect 6977 7046 6991 7098
rect 7015 7046 7029 7098
rect 7029 7046 7041 7098
rect 7041 7046 7071 7098
rect 7095 7046 7105 7098
rect 7105 7046 7151 7098
rect 6855 7044 6911 7046
rect 6935 7044 6991 7046
rect 7015 7044 7071 7046
rect 7095 7044 7151 7046
rect 10788 7098 10844 7100
rect 10868 7098 10924 7100
rect 10948 7098 11004 7100
rect 11028 7098 11084 7100
rect 10788 7046 10834 7098
rect 10834 7046 10844 7098
rect 10868 7046 10898 7098
rect 10898 7046 10910 7098
rect 10910 7046 10924 7098
rect 10948 7046 10962 7098
rect 10962 7046 10974 7098
rect 10974 7046 11004 7098
rect 11028 7046 11038 7098
rect 11038 7046 11084 7098
rect 10788 7044 10844 7046
rect 10868 7044 10924 7046
rect 10948 7044 11004 7046
rect 11028 7044 11084 7046
rect 14721 7098 14777 7100
rect 14801 7098 14857 7100
rect 14881 7098 14937 7100
rect 14961 7098 15017 7100
rect 14721 7046 14767 7098
rect 14767 7046 14777 7098
rect 14801 7046 14831 7098
rect 14831 7046 14843 7098
rect 14843 7046 14857 7098
rect 14881 7046 14895 7098
rect 14895 7046 14907 7098
rect 14907 7046 14937 7098
rect 14961 7046 14971 7098
rect 14971 7046 15017 7098
rect 14721 7044 14777 7046
rect 14801 7044 14857 7046
rect 14881 7044 14937 7046
rect 14961 7044 15017 7046
rect 4888 6554 4944 6556
rect 4968 6554 5024 6556
rect 5048 6554 5104 6556
rect 5128 6554 5184 6556
rect 4888 6502 4934 6554
rect 4934 6502 4944 6554
rect 4968 6502 4998 6554
rect 4998 6502 5010 6554
rect 5010 6502 5024 6554
rect 5048 6502 5062 6554
rect 5062 6502 5074 6554
rect 5074 6502 5104 6554
rect 5128 6502 5138 6554
rect 5138 6502 5184 6554
rect 4888 6500 4944 6502
rect 4968 6500 5024 6502
rect 5048 6500 5104 6502
rect 5128 6500 5184 6502
rect 8821 6554 8877 6556
rect 8901 6554 8957 6556
rect 8981 6554 9037 6556
rect 9061 6554 9117 6556
rect 8821 6502 8867 6554
rect 8867 6502 8877 6554
rect 8901 6502 8931 6554
rect 8931 6502 8943 6554
rect 8943 6502 8957 6554
rect 8981 6502 8995 6554
rect 8995 6502 9007 6554
rect 9007 6502 9037 6554
rect 9061 6502 9071 6554
rect 9071 6502 9117 6554
rect 8821 6500 8877 6502
rect 8901 6500 8957 6502
rect 8981 6500 9037 6502
rect 9061 6500 9117 6502
rect 12754 6554 12810 6556
rect 12834 6554 12890 6556
rect 12914 6554 12970 6556
rect 12994 6554 13050 6556
rect 12754 6502 12800 6554
rect 12800 6502 12810 6554
rect 12834 6502 12864 6554
rect 12864 6502 12876 6554
rect 12876 6502 12890 6554
rect 12914 6502 12928 6554
rect 12928 6502 12940 6554
rect 12940 6502 12970 6554
rect 12994 6502 13004 6554
rect 13004 6502 13050 6554
rect 12754 6500 12810 6502
rect 12834 6500 12890 6502
rect 12914 6500 12970 6502
rect 12994 6500 13050 6502
rect 16687 6554 16743 6556
rect 16767 6554 16823 6556
rect 16847 6554 16903 6556
rect 16927 6554 16983 6556
rect 16687 6502 16733 6554
rect 16733 6502 16743 6554
rect 16767 6502 16797 6554
rect 16797 6502 16809 6554
rect 16809 6502 16823 6554
rect 16847 6502 16861 6554
rect 16861 6502 16873 6554
rect 16873 6502 16903 6554
rect 16927 6502 16937 6554
rect 16937 6502 16983 6554
rect 16687 6500 16743 6502
rect 16767 6500 16823 6502
rect 16847 6500 16903 6502
rect 16927 6500 16983 6502
rect 2922 6010 2978 6012
rect 3002 6010 3058 6012
rect 3082 6010 3138 6012
rect 3162 6010 3218 6012
rect 2922 5958 2968 6010
rect 2968 5958 2978 6010
rect 3002 5958 3032 6010
rect 3032 5958 3044 6010
rect 3044 5958 3058 6010
rect 3082 5958 3096 6010
rect 3096 5958 3108 6010
rect 3108 5958 3138 6010
rect 3162 5958 3172 6010
rect 3172 5958 3218 6010
rect 2922 5956 2978 5958
rect 3002 5956 3058 5958
rect 3082 5956 3138 5958
rect 3162 5956 3218 5958
rect 6855 6010 6911 6012
rect 6935 6010 6991 6012
rect 7015 6010 7071 6012
rect 7095 6010 7151 6012
rect 6855 5958 6901 6010
rect 6901 5958 6911 6010
rect 6935 5958 6965 6010
rect 6965 5958 6977 6010
rect 6977 5958 6991 6010
rect 7015 5958 7029 6010
rect 7029 5958 7041 6010
rect 7041 5958 7071 6010
rect 7095 5958 7105 6010
rect 7105 5958 7151 6010
rect 6855 5956 6911 5958
rect 6935 5956 6991 5958
rect 7015 5956 7071 5958
rect 7095 5956 7151 5958
rect 10788 6010 10844 6012
rect 10868 6010 10924 6012
rect 10948 6010 11004 6012
rect 11028 6010 11084 6012
rect 10788 5958 10834 6010
rect 10834 5958 10844 6010
rect 10868 5958 10898 6010
rect 10898 5958 10910 6010
rect 10910 5958 10924 6010
rect 10948 5958 10962 6010
rect 10962 5958 10974 6010
rect 10974 5958 11004 6010
rect 11028 5958 11038 6010
rect 11038 5958 11084 6010
rect 10788 5956 10844 5958
rect 10868 5956 10924 5958
rect 10948 5956 11004 5958
rect 11028 5956 11084 5958
rect 14721 6010 14777 6012
rect 14801 6010 14857 6012
rect 14881 6010 14937 6012
rect 14961 6010 15017 6012
rect 14721 5958 14767 6010
rect 14767 5958 14777 6010
rect 14801 5958 14831 6010
rect 14831 5958 14843 6010
rect 14843 5958 14857 6010
rect 14881 5958 14895 6010
rect 14895 5958 14907 6010
rect 14907 5958 14937 6010
rect 14961 5958 14971 6010
rect 14971 5958 15017 6010
rect 14721 5956 14777 5958
rect 14801 5956 14857 5958
rect 14881 5956 14937 5958
rect 14961 5956 15017 5958
rect 4888 5466 4944 5468
rect 4968 5466 5024 5468
rect 5048 5466 5104 5468
rect 5128 5466 5184 5468
rect 4888 5414 4934 5466
rect 4934 5414 4944 5466
rect 4968 5414 4998 5466
rect 4998 5414 5010 5466
rect 5010 5414 5024 5466
rect 5048 5414 5062 5466
rect 5062 5414 5074 5466
rect 5074 5414 5104 5466
rect 5128 5414 5138 5466
rect 5138 5414 5184 5466
rect 4888 5412 4944 5414
rect 4968 5412 5024 5414
rect 5048 5412 5104 5414
rect 5128 5412 5184 5414
rect 8821 5466 8877 5468
rect 8901 5466 8957 5468
rect 8981 5466 9037 5468
rect 9061 5466 9117 5468
rect 8821 5414 8867 5466
rect 8867 5414 8877 5466
rect 8901 5414 8931 5466
rect 8931 5414 8943 5466
rect 8943 5414 8957 5466
rect 8981 5414 8995 5466
rect 8995 5414 9007 5466
rect 9007 5414 9037 5466
rect 9061 5414 9071 5466
rect 9071 5414 9117 5466
rect 8821 5412 8877 5414
rect 8901 5412 8957 5414
rect 8981 5412 9037 5414
rect 9061 5412 9117 5414
rect 12754 5466 12810 5468
rect 12834 5466 12890 5468
rect 12914 5466 12970 5468
rect 12994 5466 13050 5468
rect 12754 5414 12800 5466
rect 12800 5414 12810 5466
rect 12834 5414 12864 5466
rect 12864 5414 12876 5466
rect 12876 5414 12890 5466
rect 12914 5414 12928 5466
rect 12928 5414 12940 5466
rect 12940 5414 12970 5466
rect 12994 5414 13004 5466
rect 13004 5414 13050 5466
rect 12754 5412 12810 5414
rect 12834 5412 12890 5414
rect 12914 5412 12970 5414
rect 12994 5412 13050 5414
rect 16687 5466 16743 5468
rect 16767 5466 16823 5468
rect 16847 5466 16903 5468
rect 16927 5466 16983 5468
rect 16687 5414 16733 5466
rect 16733 5414 16743 5466
rect 16767 5414 16797 5466
rect 16797 5414 16809 5466
rect 16809 5414 16823 5466
rect 16847 5414 16861 5466
rect 16861 5414 16873 5466
rect 16873 5414 16903 5466
rect 16927 5414 16937 5466
rect 16937 5414 16983 5466
rect 16687 5412 16743 5414
rect 16767 5412 16823 5414
rect 16847 5412 16903 5414
rect 16927 5412 16983 5414
rect 2922 4922 2978 4924
rect 3002 4922 3058 4924
rect 3082 4922 3138 4924
rect 3162 4922 3218 4924
rect 2922 4870 2968 4922
rect 2968 4870 2978 4922
rect 3002 4870 3032 4922
rect 3032 4870 3044 4922
rect 3044 4870 3058 4922
rect 3082 4870 3096 4922
rect 3096 4870 3108 4922
rect 3108 4870 3138 4922
rect 3162 4870 3172 4922
rect 3172 4870 3218 4922
rect 2922 4868 2978 4870
rect 3002 4868 3058 4870
rect 3082 4868 3138 4870
rect 3162 4868 3218 4870
rect 6855 4922 6911 4924
rect 6935 4922 6991 4924
rect 7015 4922 7071 4924
rect 7095 4922 7151 4924
rect 6855 4870 6901 4922
rect 6901 4870 6911 4922
rect 6935 4870 6965 4922
rect 6965 4870 6977 4922
rect 6977 4870 6991 4922
rect 7015 4870 7029 4922
rect 7029 4870 7041 4922
rect 7041 4870 7071 4922
rect 7095 4870 7105 4922
rect 7105 4870 7151 4922
rect 6855 4868 6911 4870
rect 6935 4868 6991 4870
rect 7015 4868 7071 4870
rect 7095 4868 7151 4870
rect 10788 4922 10844 4924
rect 10868 4922 10924 4924
rect 10948 4922 11004 4924
rect 11028 4922 11084 4924
rect 10788 4870 10834 4922
rect 10834 4870 10844 4922
rect 10868 4870 10898 4922
rect 10898 4870 10910 4922
rect 10910 4870 10924 4922
rect 10948 4870 10962 4922
rect 10962 4870 10974 4922
rect 10974 4870 11004 4922
rect 11028 4870 11038 4922
rect 11038 4870 11084 4922
rect 10788 4868 10844 4870
rect 10868 4868 10924 4870
rect 10948 4868 11004 4870
rect 11028 4868 11084 4870
rect 14721 4922 14777 4924
rect 14801 4922 14857 4924
rect 14881 4922 14937 4924
rect 14961 4922 15017 4924
rect 14721 4870 14767 4922
rect 14767 4870 14777 4922
rect 14801 4870 14831 4922
rect 14831 4870 14843 4922
rect 14843 4870 14857 4922
rect 14881 4870 14895 4922
rect 14895 4870 14907 4922
rect 14907 4870 14937 4922
rect 14961 4870 14971 4922
rect 14971 4870 15017 4922
rect 14721 4868 14777 4870
rect 14801 4868 14857 4870
rect 14881 4868 14937 4870
rect 14961 4868 15017 4870
rect 4888 4378 4944 4380
rect 4968 4378 5024 4380
rect 5048 4378 5104 4380
rect 5128 4378 5184 4380
rect 4888 4326 4934 4378
rect 4934 4326 4944 4378
rect 4968 4326 4998 4378
rect 4998 4326 5010 4378
rect 5010 4326 5024 4378
rect 5048 4326 5062 4378
rect 5062 4326 5074 4378
rect 5074 4326 5104 4378
rect 5128 4326 5138 4378
rect 5138 4326 5184 4378
rect 4888 4324 4944 4326
rect 4968 4324 5024 4326
rect 5048 4324 5104 4326
rect 5128 4324 5184 4326
rect 8821 4378 8877 4380
rect 8901 4378 8957 4380
rect 8981 4378 9037 4380
rect 9061 4378 9117 4380
rect 8821 4326 8867 4378
rect 8867 4326 8877 4378
rect 8901 4326 8931 4378
rect 8931 4326 8943 4378
rect 8943 4326 8957 4378
rect 8981 4326 8995 4378
rect 8995 4326 9007 4378
rect 9007 4326 9037 4378
rect 9061 4326 9071 4378
rect 9071 4326 9117 4378
rect 8821 4324 8877 4326
rect 8901 4324 8957 4326
rect 8981 4324 9037 4326
rect 9061 4324 9117 4326
rect 12754 4378 12810 4380
rect 12834 4378 12890 4380
rect 12914 4378 12970 4380
rect 12994 4378 13050 4380
rect 12754 4326 12800 4378
rect 12800 4326 12810 4378
rect 12834 4326 12864 4378
rect 12864 4326 12876 4378
rect 12876 4326 12890 4378
rect 12914 4326 12928 4378
rect 12928 4326 12940 4378
rect 12940 4326 12970 4378
rect 12994 4326 13004 4378
rect 13004 4326 13050 4378
rect 12754 4324 12810 4326
rect 12834 4324 12890 4326
rect 12914 4324 12970 4326
rect 12994 4324 13050 4326
rect 16687 4378 16743 4380
rect 16767 4378 16823 4380
rect 16847 4378 16903 4380
rect 16927 4378 16983 4380
rect 16687 4326 16733 4378
rect 16733 4326 16743 4378
rect 16767 4326 16797 4378
rect 16797 4326 16809 4378
rect 16809 4326 16823 4378
rect 16847 4326 16861 4378
rect 16861 4326 16873 4378
rect 16873 4326 16903 4378
rect 16927 4326 16937 4378
rect 16937 4326 16983 4378
rect 16687 4324 16743 4326
rect 16767 4324 16823 4326
rect 16847 4324 16903 4326
rect 16927 4324 16983 4326
rect 2922 3834 2978 3836
rect 3002 3834 3058 3836
rect 3082 3834 3138 3836
rect 3162 3834 3218 3836
rect 2922 3782 2968 3834
rect 2968 3782 2978 3834
rect 3002 3782 3032 3834
rect 3032 3782 3044 3834
rect 3044 3782 3058 3834
rect 3082 3782 3096 3834
rect 3096 3782 3108 3834
rect 3108 3782 3138 3834
rect 3162 3782 3172 3834
rect 3172 3782 3218 3834
rect 2922 3780 2978 3782
rect 3002 3780 3058 3782
rect 3082 3780 3138 3782
rect 3162 3780 3218 3782
rect 6855 3834 6911 3836
rect 6935 3834 6991 3836
rect 7015 3834 7071 3836
rect 7095 3834 7151 3836
rect 6855 3782 6901 3834
rect 6901 3782 6911 3834
rect 6935 3782 6965 3834
rect 6965 3782 6977 3834
rect 6977 3782 6991 3834
rect 7015 3782 7029 3834
rect 7029 3782 7041 3834
rect 7041 3782 7071 3834
rect 7095 3782 7105 3834
rect 7105 3782 7151 3834
rect 6855 3780 6911 3782
rect 6935 3780 6991 3782
rect 7015 3780 7071 3782
rect 7095 3780 7151 3782
rect 10788 3834 10844 3836
rect 10868 3834 10924 3836
rect 10948 3834 11004 3836
rect 11028 3834 11084 3836
rect 10788 3782 10834 3834
rect 10834 3782 10844 3834
rect 10868 3782 10898 3834
rect 10898 3782 10910 3834
rect 10910 3782 10924 3834
rect 10948 3782 10962 3834
rect 10962 3782 10974 3834
rect 10974 3782 11004 3834
rect 11028 3782 11038 3834
rect 11038 3782 11084 3834
rect 10788 3780 10844 3782
rect 10868 3780 10924 3782
rect 10948 3780 11004 3782
rect 11028 3780 11084 3782
rect 14721 3834 14777 3836
rect 14801 3834 14857 3836
rect 14881 3834 14937 3836
rect 14961 3834 15017 3836
rect 14721 3782 14767 3834
rect 14767 3782 14777 3834
rect 14801 3782 14831 3834
rect 14831 3782 14843 3834
rect 14843 3782 14857 3834
rect 14881 3782 14895 3834
rect 14895 3782 14907 3834
rect 14907 3782 14937 3834
rect 14961 3782 14971 3834
rect 14971 3782 15017 3834
rect 14721 3780 14777 3782
rect 14801 3780 14857 3782
rect 14881 3780 14937 3782
rect 14961 3780 15017 3782
rect 4888 3290 4944 3292
rect 4968 3290 5024 3292
rect 5048 3290 5104 3292
rect 5128 3290 5184 3292
rect 4888 3238 4934 3290
rect 4934 3238 4944 3290
rect 4968 3238 4998 3290
rect 4998 3238 5010 3290
rect 5010 3238 5024 3290
rect 5048 3238 5062 3290
rect 5062 3238 5074 3290
rect 5074 3238 5104 3290
rect 5128 3238 5138 3290
rect 5138 3238 5184 3290
rect 4888 3236 4944 3238
rect 4968 3236 5024 3238
rect 5048 3236 5104 3238
rect 5128 3236 5184 3238
rect 8821 3290 8877 3292
rect 8901 3290 8957 3292
rect 8981 3290 9037 3292
rect 9061 3290 9117 3292
rect 8821 3238 8867 3290
rect 8867 3238 8877 3290
rect 8901 3238 8931 3290
rect 8931 3238 8943 3290
rect 8943 3238 8957 3290
rect 8981 3238 8995 3290
rect 8995 3238 9007 3290
rect 9007 3238 9037 3290
rect 9061 3238 9071 3290
rect 9071 3238 9117 3290
rect 8821 3236 8877 3238
rect 8901 3236 8957 3238
rect 8981 3236 9037 3238
rect 9061 3236 9117 3238
rect 12754 3290 12810 3292
rect 12834 3290 12890 3292
rect 12914 3290 12970 3292
rect 12994 3290 13050 3292
rect 12754 3238 12800 3290
rect 12800 3238 12810 3290
rect 12834 3238 12864 3290
rect 12864 3238 12876 3290
rect 12876 3238 12890 3290
rect 12914 3238 12928 3290
rect 12928 3238 12940 3290
rect 12940 3238 12970 3290
rect 12994 3238 13004 3290
rect 13004 3238 13050 3290
rect 12754 3236 12810 3238
rect 12834 3236 12890 3238
rect 12914 3236 12970 3238
rect 12994 3236 13050 3238
rect 16687 3290 16743 3292
rect 16767 3290 16823 3292
rect 16847 3290 16903 3292
rect 16927 3290 16983 3292
rect 16687 3238 16733 3290
rect 16733 3238 16743 3290
rect 16767 3238 16797 3290
rect 16797 3238 16809 3290
rect 16809 3238 16823 3290
rect 16847 3238 16861 3290
rect 16861 3238 16873 3290
rect 16873 3238 16903 3290
rect 16927 3238 16937 3290
rect 16937 3238 16983 3290
rect 16687 3236 16743 3238
rect 16767 3236 16823 3238
rect 16847 3236 16903 3238
rect 16927 3236 16983 3238
rect 2922 2746 2978 2748
rect 3002 2746 3058 2748
rect 3082 2746 3138 2748
rect 3162 2746 3218 2748
rect 2922 2694 2968 2746
rect 2968 2694 2978 2746
rect 3002 2694 3032 2746
rect 3032 2694 3044 2746
rect 3044 2694 3058 2746
rect 3082 2694 3096 2746
rect 3096 2694 3108 2746
rect 3108 2694 3138 2746
rect 3162 2694 3172 2746
rect 3172 2694 3218 2746
rect 2922 2692 2978 2694
rect 3002 2692 3058 2694
rect 3082 2692 3138 2694
rect 3162 2692 3218 2694
rect 6855 2746 6911 2748
rect 6935 2746 6991 2748
rect 7015 2746 7071 2748
rect 7095 2746 7151 2748
rect 6855 2694 6901 2746
rect 6901 2694 6911 2746
rect 6935 2694 6965 2746
rect 6965 2694 6977 2746
rect 6977 2694 6991 2746
rect 7015 2694 7029 2746
rect 7029 2694 7041 2746
rect 7041 2694 7071 2746
rect 7095 2694 7105 2746
rect 7105 2694 7151 2746
rect 6855 2692 6911 2694
rect 6935 2692 6991 2694
rect 7015 2692 7071 2694
rect 7095 2692 7151 2694
rect 10788 2746 10844 2748
rect 10868 2746 10924 2748
rect 10948 2746 11004 2748
rect 11028 2746 11084 2748
rect 10788 2694 10834 2746
rect 10834 2694 10844 2746
rect 10868 2694 10898 2746
rect 10898 2694 10910 2746
rect 10910 2694 10924 2746
rect 10948 2694 10962 2746
rect 10962 2694 10974 2746
rect 10974 2694 11004 2746
rect 11028 2694 11038 2746
rect 11038 2694 11084 2746
rect 10788 2692 10844 2694
rect 10868 2692 10924 2694
rect 10948 2692 11004 2694
rect 11028 2692 11084 2694
rect 14721 2746 14777 2748
rect 14801 2746 14857 2748
rect 14881 2746 14937 2748
rect 14961 2746 15017 2748
rect 14721 2694 14767 2746
rect 14767 2694 14777 2746
rect 14801 2694 14831 2746
rect 14831 2694 14843 2746
rect 14843 2694 14857 2746
rect 14881 2694 14895 2746
rect 14895 2694 14907 2746
rect 14907 2694 14937 2746
rect 14961 2694 14971 2746
rect 14971 2694 15017 2746
rect 14721 2692 14777 2694
rect 14801 2692 14857 2694
rect 14881 2692 14937 2694
rect 14961 2692 15017 2694
rect 1766 2252 1768 2272
rect 1768 2252 1820 2272
rect 1820 2252 1822 2272
rect 1766 2216 1822 2252
rect 4888 2202 4944 2204
rect 4968 2202 5024 2204
rect 5048 2202 5104 2204
rect 5128 2202 5184 2204
rect 4888 2150 4934 2202
rect 4934 2150 4944 2202
rect 4968 2150 4998 2202
rect 4998 2150 5010 2202
rect 5010 2150 5024 2202
rect 5048 2150 5062 2202
rect 5062 2150 5074 2202
rect 5074 2150 5104 2202
rect 5128 2150 5138 2202
rect 5138 2150 5184 2202
rect 4888 2148 4944 2150
rect 4968 2148 5024 2150
rect 5048 2148 5104 2150
rect 5128 2148 5184 2150
rect 8821 2202 8877 2204
rect 8901 2202 8957 2204
rect 8981 2202 9037 2204
rect 9061 2202 9117 2204
rect 8821 2150 8867 2202
rect 8867 2150 8877 2202
rect 8901 2150 8931 2202
rect 8931 2150 8943 2202
rect 8943 2150 8957 2202
rect 8981 2150 8995 2202
rect 8995 2150 9007 2202
rect 9007 2150 9037 2202
rect 9061 2150 9071 2202
rect 9071 2150 9117 2202
rect 8821 2148 8877 2150
rect 8901 2148 8957 2150
rect 8981 2148 9037 2150
rect 9061 2148 9117 2150
rect 12754 2202 12810 2204
rect 12834 2202 12890 2204
rect 12914 2202 12970 2204
rect 12994 2202 13050 2204
rect 12754 2150 12800 2202
rect 12800 2150 12810 2202
rect 12834 2150 12864 2202
rect 12864 2150 12876 2202
rect 12876 2150 12890 2202
rect 12914 2150 12928 2202
rect 12928 2150 12940 2202
rect 12940 2150 12970 2202
rect 12994 2150 13004 2202
rect 13004 2150 13050 2202
rect 12754 2148 12810 2150
rect 12834 2148 12890 2150
rect 12914 2148 12970 2150
rect 12994 2148 13050 2150
rect 16687 2202 16743 2204
rect 16767 2202 16823 2204
rect 16847 2202 16903 2204
rect 16927 2202 16983 2204
rect 16687 2150 16733 2202
rect 16733 2150 16743 2202
rect 16767 2150 16797 2202
rect 16797 2150 16809 2202
rect 16809 2150 16823 2202
rect 16847 2150 16861 2202
rect 16861 2150 16873 2202
rect 16873 2150 16903 2202
rect 16927 2150 16937 2202
rect 16937 2150 16983 2202
rect 16687 2148 16743 2150
rect 16767 2148 16823 2150
rect 16847 2148 16903 2150
rect 16927 2148 16983 2150
<< metal3 >>
rect 2912 15808 3228 15809
rect 0 15738 800 15768
rect 2912 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3228 15808
rect 2912 15743 3228 15744
rect 6845 15808 7161 15809
rect 6845 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7161 15808
rect 6845 15743 7161 15744
rect 10778 15808 11094 15809
rect 10778 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11094 15808
rect 10778 15743 11094 15744
rect 14711 15808 15027 15809
rect 14711 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15027 15808
rect 14711 15743 15027 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15648 800 15678
rect 2773 15675 2839 15678
rect 4878 15264 5194 15265
rect 4878 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5194 15264
rect 4878 15199 5194 15200
rect 8811 15264 9127 15265
rect 8811 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9127 15264
rect 8811 15199 9127 15200
rect 12744 15264 13060 15265
rect 12744 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13060 15264
rect 12744 15199 13060 15200
rect 16677 15264 16993 15265
rect 16677 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16993 15264
rect 16677 15199 16993 15200
rect 5717 15058 5783 15061
rect 6545 15058 6611 15061
rect 5717 15056 6611 15058
rect 5717 15000 5722 15056
rect 5778 15000 6550 15056
rect 6606 15000 6611 15056
rect 5717 14998 6611 15000
rect 5717 14995 5783 14998
rect 6545 14995 6611 14998
rect 2912 14720 3228 14721
rect 2912 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3228 14720
rect 2912 14655 3228 14656
rect 6845 14720 7161 14721
rect 6845 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7161 14720
rect 6845 14655 7161 14656
rect 10778 14720 11094 14721
rect 10778 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11094 14720
rect 10778 14655 11094 14656
rect 14711 14720 15027 14721
rect 14711 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15027 14720
rect 14711 14655 15027 14656
rect 4878 14176 5194 14177
rect 4878 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5194 14176
rect 4878 14111 5194 14112
rect 8811 14176 9127 14177
rect 8811 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9127 14176
rect 8811 14111 9127 14112
rect 12744 14176 13060 14177
rect 12744 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13060 14176
rect 12744 14111 13060 14112
rect 16677 14176 16993 14177
rect 16677 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16993 14176
rect 16677 14111 16993 14112
rect 2221 13970 2287 13973
rect 4061 13970 4127 13973
rect 5625 13970 5691 13973
rect 7833 13970 7899 13973
rect 2221 13968 7899 13970
rect 2221 13912 2226 13968
rect 2282 13912 4066 13968
rect 4122 13912 5630 13968
rect 5686 13912 7838 13968
rect 7894 13912 7899 13968
rect 2221 13910 7899 13912
rect 2221 13907 2287 13910
rect 4061 13907 4127 13910
rect 5625 13907 5691 13910
rect 7833 13907 7899 13910
rect 2912 13632 3228 13633
rect 2912 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3228 13632
rect 2912 13567 3228 13568
rect 6845 13632 7161 13633
rect 6845 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7161 13632
rect 6845 13567 7161 13568
rect 10778 13632 11094 13633
rect 10778 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11094 13632
rect 10778 13567 11094 13568
rect 14711 13632 15027 13633
rect 14711 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15027 13632
rect 14711 13567 15027 13568
rect 4878 13088 5194 13089
rect 4878 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5194 13088
rect 4878 13023 5194 13024
rect 8811 13088 9127 13089
rect 8811 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9127 13088
rect 8811 13023 9127 13024
rect 12744 13088 13060 13089
rect 12744 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13060 13088
rect 12744 13023 13060 13024
rect 16677 13088 16993 13089
rect 16677 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16993 13088
rect 16677 13023 16993 13024
rect 2912 12544 3228 12545
rect 2912 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3228 12544
rect 2912 12479 3228 12480
rect 6845 12544 7161 12545
rect 6845 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7161 12544
rect 6845 12479 7161 12480
rect 10778 12544 11094 12545
rect 10778 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11094 12544
rect 10778 12479 11094 12480
rect 14711 12544 15027 12545
rect 14711 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15027 12544
rect 14711 12479 15027 12480
rect 4878 12000 5194 12001
rect 4878 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5194 12000
rect 4878 11935 5194 11936
rect 8811 12000 9127 12001
rect 8811 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9127 12000
rect 8811 11935 9127 11936
rect 12744 12000 13060 12001
rect 12744 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13060 12000
rect 12744 11935 13060 11936
rect 16677 12000 16993 12001
rect 16677 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16993 12000
rect 16677 11935 16993 11936
rect 2912 11456 3228 11457
rect 2912 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3228 11456
rect 2912 11391 3228 11392
rect 6845 11456 7161 11457
rect 6845 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7161 11456
rect 6845 11391 7161 11392
rect 10778 11456 11094 11457
rect 10778 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11094 11456
rect 10778 11391 11094 11392
rect 14711 11456 15027 11457
rect 14711 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15027 11456
rect 14711 11391 15027 11392
rect 0 11250 800 11280
rect 1669 11250 1735 11253
rect 0 11248 1735 11250
rect 0 11192 1674 11248
rect 1730 11192 1735 11248
rect 0 11190 1735 11192
rect 0 11160 800 11190
rect 1669 11187 1735 11190
rect 4878 10912 5194 10913
rect 4878 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5194 10912
rect 4878 10847 5194 10848
rect 8811 10912 9127 10913
rect 8811 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9127 10912
rect 8811 10847 9127 10848
rect 12744 10912 13060 10913
rect 12744 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13060 10912
rect 12744 10847 13060 10848
rect 16677 10912 16993 10913
rect 16677 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16993 10912
rect 16677 10847 16993 10848
rect 2912 10368 3228 10369
rect 2912 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3228 10368
rect 2912 10303 3228 10304
rect 6845 10368 7161 10369
rect 6845 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7161 10368
rect 6845 10303 7161 10304
rect 10778 10368 11094 10369
rect 10778 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11094 10368
rect 10778 10303 11094 10304
rect 14711 10368 15027 10369
rect 14711 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15027 10368
rect 14711 10303 15027 10304
rect 4878 9824 5194 9825
rect 4878 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5194 9824
rect 4878 9759 5194 9760
rect 8811 9824 9127 9825
rect 8811 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9127 9824
rect 8811 9759 9127 9760
rect 12744 9824 13060 9825
rect 12744 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13060 9824
rect 12744 9759 13060 9760
rect 16677 9824 16993 9825
rect 16677 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16993 9824
rect 16677 9759 16993 9760
rect 2912 9280 3228 9281
rect 2912 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3228 9280
rect 2912 9215 3228 9216
rect 6845 9280 7161 9281
rect 6845 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7161 9280
rect 6845 9215 7161 9216
rect 10778 9280 11094 9281
rect 10778 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11094 9280
rect 10778 9215 11094 9216
rect 14711 9280 15027 9281
rect 14711 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15027 9280
rect 14711 9215 15027 9216
rect 4878 8736 5194 8737
rect 4878 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5194 8736
rect 4878 8671 5194 8672
rect 8811 8736 9127 8737
rect 8811 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9127 8736
rect 8811 8671 9127 8672
rect 12744 8736 13060 8737
rect 12744 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13060 8736
rect 12744 8671 13060 8672
rect 16677 8736 16993 8737
rect 16677 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16993 8736
rect 16677 8671 16993 8672
rect 2912 8192 3228 8193
rect 2912 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3228 8192
rect 2912 8127 3228 8128
rect 6845 8192 7161 8193
rect 6845 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7161 8192
rect 6845 8127 7161 8128
rect 10778 8192 11094 8193
rect 10778 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11094 8192
rect 10778 8127 11094 8128
rect 14711 8192 15027 8193
rect 14711 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15027 8192
rect 14711 8127 15027 8128
rect 4878 7648 5194 7649
rect 4878 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5194 7648
rect 4878 7583 5194 7584
rect 8811 7648 9127 7649
rect 8811 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9127 7648
rect 8811 7583 9127 7584
rect 12744 7648 13060 7649
rect 12744 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13060 7648
rect 12744 7583 13060 7584
rect 16677 7648 16993 7649
rect 16677 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16993 7648
rect 16677 7583 16993 7584
rect 2912 7104 3228 7105
rect 2912 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3228 7104
rect 2912 7039 3228 7040
rect 6845 7104 7161 7105
rect 6845 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7161 7104
rect 6845 7039 7161 7040
rect 10778 7104 11094 7105
rect 10778 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11094 7104
rect 10778 7039 11094 7040
rect 14711 7104 15027 7105
rect 14711 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15027 7104
rect 14711 7039 15027 7040
rect 0 6762 800 6792
rect 1485 6762 1551 6765
rect 0 6760 1551 6762
rect 0 6704 1490 6760
rect 1546 6704 1551 6760
rect 0 6702 1551 6704
rect 0 6672 800 6702
rect 1485 6699 1551 6702
rect 4878 6560 5194 6561
rect 4878 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5194 6560
rect 4878 6495 5194 6496
rect 8811 6560 9127 6561
rect 8811 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9127 6560
rect 8811 6495 9127 6496
rect 12744 6560 13060 6561
rect 12744 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13060 6560
rect 12744 6495 13060 6496
rect 16677 6560 16993 6561
rect 16677 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16993 6560
rect 16677 6495 16993 6496
rect 2912 6016 3228 6017
rect 2912 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3228 6016
rect 2912 5951 3228 5952
rect 6845 6016 7161 6017
rect 6845 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7161 6016
rect 6845 5951 7161 5952
rect 10778 6016 11094 6017
rect 10778 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11094 6016
rect 10778 5951 11094 5952
rect 14711 6016 15027 6017
rect 14711 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15027 6016
rect 14711 5951 15027 5952
rect 4878 5472 5194 5473
rect 4878 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5194 5472
rect 4878 5407 5194 5408
rect 8811 5472 9127 5473
rect 8811 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9127 5472
rect 8811 5407 9127 5408
rect 12744 5472 13060 5473
rect 12744 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13060 5472
rect 12744 5407 13060 5408
rect 16677 5472 16993 5473
rect 16677 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16993 5472
rect 16677 5407 16993 5408
rect 2912 4928 3228 4929
rect 2912 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3228 4928
rect 2912 4863 3228 4864
rect 6845 4928 7161 4929
rect 6845 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7161 4928
rect 6845 4863 7161 4864
rect 10778 4928 11094 4929
rect 10778 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11094 4928
rect 10778 4863 11094 4864
rect 14711 4928 15027 4929
rect 14711 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15027 4928
rect 14711 4863 15027 4864
rect 4878 4384 5194 4385
rect 4878 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5194 4384
rect 4878 4319 5194 4320
rect 8811 4384 9127 4385
rect 8811 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9127 4384
rect 8811 4319 9127 4320
rect 12744 4384 13060 4385
rect 12744 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13060 4384
rect 12744 4319 13060 4320
rect 16677 4384 16993 4385
rect 16677 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16993 4384
rect 16677 4319 16993 4320
rect 2912 3840 3228 3841
rect 2912 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3228 3840
rect 2912 3775 3228 3776
rect 6845 3840 7161 3841
rect 6845 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7161 3840
rect 6845 3775 7161 3776
rect 10778 3840 11094 3841
rect 10778 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11094 3840
rect 10778 3775 11094 3776
rect 14711 3840 15027 3841
rect 14711 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15027 3840
rect 14711 3775 15027 3776
rect 4878 3296 5194 3297
rect 4878 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5194 3296
rect 4878 3231 5194 3232
rect 8811 3296 9127 3297
rect 8811 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9127 3296
rect 8811 3231 9127 3232
rect 12744 3296 13060 3297
rect 12744 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13060 3296
rect 12744 3231 13060 3232
rect 16677 3296 16993 3297
rect 16677 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16993 3296
rect 16677 3231 16993 3232
rect 2912 2752 3228 2753
rect 2912 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3228 2752
rect 2912 2687 3228 2688
rect 6845 2752 7161 2753
rect 6845 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7161 2752
rect 6845 2687 7161 2688
rect 10778 2752 11094 2753
rect 10778 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11094 2752
rect 10778 2687 11094 2688
rect 14711 2752 15027 2753
rect 14711 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15027 2752
rect 14711 2687 15027 2688
rect 0 2274 800 2304
rect 1761 2274 1827 2277
rect 0 2272 1827 2274
rect 0 2216 1766 2272
rect 1822 2216 1827 2272
rect 0 2214 1827 2216
rect 0 2184 800 2214
rect 1761 2211 1827 2214
rect 4878 2208 5194 2209
rect 4878 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5194 2208
rect 4878 2143 5194 2144
rect 8811 2208 9127 2209
rect 8811 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9127 2208
rect 8811 2143 9127 2144
rect 12744 2208 13060 2209
rect 12744 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13060 2208
rect 12744 2143 13060 2144
rect 16677 2208 16993 2209
rect 16677 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16993 2208
rect 16677 2143 16993 2144
<< via3 >>
rect 2918 15804 2982 15808
rect 2918 15748 2922 15804
rect 2922 15748 2978 15804
rect 2978 15748 2982 15804
rect 2918 15744 2982 15748
rect 2998 15804 3062 15808
rect 2998 15748 3002 15804
rect 3002 15748 3058 15804
rect 3058 15748 3062 15804
rect 2998 15744 3062 15748
rect 3078 15804 3142 15808
rect 3078 15748 3082 15804
rect 3082 15748 3138 15804
rect 3138 15748 3142 15804
rect 3078 15744 3142 15748
rect 3158 15804 3222 15808
rect 3158 15748 3162 15804
rect 3162 15748 3218 15804
rect 3218 15748 3222 15804
rect 3158 15744 3222 15748
rect 6851 15804 6915 15808
rect 6851 15748 6855 15804
rect 6855 15748 6911 15804
rect 6911 15748 6915 15804
rect 6851 15744 6915 15748
rect 6931 15804 6995 15808
rect 6931 15748 6935 15804
rect 6935 15748 6991 15804
rect 6991 15748 6995 15804
rect 6931 15744 6995 15748
rect 7011 15804 7075 15808
rect 7011 15748 7015 15804
rect 7015 15748 7071 15804
rect 7071 15748 7075 15804
rect 7011 15744 7075 15748
rect 7091 15804 7155 15808
rect 7091 15748 7095 15804
rect 7095 15748 7151 15804
rect 7151 15748 7155 15804
rect 7091 15744 7155 15748
rect 10784 15804 10848 15808
rect 10784 15748 10788 15804
rect 10788 15748 10844 15804
rect 10844 15748 10848 15804
rect 10784 15744 10848 15748
rect 10864 15804 10928 15808
rect 10864 15748 10868 15804
rect 10868 15748 10924 15804
rect 10924 15748 10928 15804
rect 10864 15744 10928 15748
rect 10944 15804 11008 15808
rect 10944 15748 10948 15804
rect 10948 15748 11004 15804
rect 11004 15748 11008 15804
rect 10944 15744 11008 15748
rect 11024 15804 11088 15808
rect 11024 15748 11028 15804
rect 11028 15748 11084 15804
rect 11084 15748 11088 15804
rect 11024 15744 11088 15748
rect 14717 15804 14781 15808
rect 14717 15748 14721 15804
rect 14721 15748 14777 15804
rect 14777 15748 14781 15804
rect 14717 15744 14781 15748
rect 14797 15804 14861 15808
rect 14797 15748 14801 15804
rect 14801 15748 14857 15804
rect 14857 15748 14861 15804
rect 14797 15744 14861 15748
rect 14877 15804 14941 15808
rect 14877 15748 14881 15804
rect 14881 15748 14937 15804
rect 14937 15748 14941 15804
rect 14877 15744 14941 15748
rect 14957 15804 15021 15808
rect 14957 15748 14961 15804
rect 14961 15748 15017 15804
rect 15017 15748 15021 15804
rect 14957 15744 15021 15748
rect 4884 15260 4948 15264
rect 4884 15204 4888 15260
rect 4888 15204 4944 15260
rect 4944 15204 4948 15260
rect 4884 15200 4948 15204
rect 4964 15260 5028 15264
rect 4964 15204 4968 15260
rect 4968 15204 5024 15260
rect 5024 15204 5028 15260
rect 4964 15200 5028 15204
rect 5044 15260 5108 15264
rect 5044 15204 5048 15260
rect 5048 15204 5104 15260
rect 5104 15204 5108 15260
rect 5044 15200 5108 15204
rect 5124 15260 5188 15264
rect 5124 15204 5128 15260
rect 5128 15204 5184 15260
rect 5184 15204 5188 15260
rect 5124 15200 5188 15204
rect 8817 15260 8881 15264
rect 8817 15204 8821 15260
rect 8821 15204 8877 15260
rect 8877 15204 8881 15260
rect 8817 15200 8881 15204
rect 8897 15260 8961 15264
rect 8897 15204 8901 15260
rect 8901 15204 8957 15260
rect 8957 15204 8961 15260
rect 8897 15200 8961 15204
rect 8977 15260 9041 15264
rect 8977 15204 8981 15260
rect 8981 15204 9037 15260
rect 9037 15204 9041 15260
rect 8977 15200 9041 15204
rect 9057 15260 9121 15264
rect 9057 15204 9061 15260
rect 9061 15204 9117 15260
rect 9117 15204 9121 15260
rect 9057 15200 9121 15204
rect 12750 15260 12814 15264
rect 12750 15204 12754 15260
rect 12754 15204 12810 15260
rect 12810 15204 12814 15260
rect 12750 15200 12814 15204
rect 12830 15260 12894 15264
rect 12830 15204 12834 15260
rect 12834 15204 12890 15260
rect 12890 15204 12894 15260
rect 12830 15200 12894 15204
rect 12910 15260 12974 15264
rect 12910 15204 12914 15260
rect 12914 15204 12970 15260
rect 12970 15204 12974 15260
rect 12910 15200 12974 15204
rect 12990 15260 13054 15264
rect 12990 15204 12994 15260
rect 12994 15204 13050 15260
rect 13050 15204 13054 15260
rect 12990 15200 13054 15204
rect 16683 15260 16747 15264
rect 16683 15204 16687 15260
rect 16687 15204 16743 15260
rect 16743 15204 16747 15260
rect 16683 15200 16747 15204
rect 16763 15260 16827 15264
rect 16763 15204 16767 15260
rect 16767 15204 16823 15260
rect 16823 15204 16827 15260
rect 16763 15200 16827 15204
rect 16843 15260 16907 15264
rect 16843 15204 16847 15260
rect 16847 15204 16903 15260
rect 16903 15204 16907 15260
rect 16843 15200 16907 15204
rect 16923 15260 16987 15264
rect 16923 15204 16927 15260
rect 16927 15204 16983 15260
rect 16983 15204 16987 15260
rect 16923 15200 16987 15204
rect 2918 14716 2982 14720
rect 2918 14660 2922 14716
rect 2922 14660 2978 14716
rect 2978 14660 2982 14716
rect 2918 14656 2982 14660
rect 2998 14716 3062 14720
rect 2998 14660 3002 14716
rect 3002 14660 3058 14716
rect 3058 14660 3062 14716
rect 2998 14656 3062 14660
rect 3078 14716 3142 14720
rect 3078 14660 3082 14716
rect 3082 14660 3138 14716
rect 3138 14660 3142 14716
rect 3078 14656 3142 14660
rect 3158 14716 3222 14720
rect 3158 14660 3162 14716
rect 3162 14660 3218 14716
rect 3218 14660 3222 14716
rect 3158 14656 3222 14660
rect 6851 14716 6915 14720
rect 6851 14660 6855 14716
rect 6855 14660 6911 14716
rect 6911 14660 6915 14716
rect 6851 14656 6915 14660
rect 6931 14716 6995 14720
rect 6931 14660 6935 14716
rect 6935 14660 6991 14716
rect 6991 14660 6995 14716
rect 6931 14656 6995 14660
rect 7011 14716 7075 14720
rect 7011 14660 7015 14716
rect 7015 14660 7071 14716
rect 7071 14660 7075 14716
rect 7011 14656 7075 14660
rect 7091 14716 7155 14720
rect 7091 14660 7095 14716
rect 7095 14660 7151 14716
rect 7151 14660 7155 14716
rect 7091 14656 7155 14660
rect 10784 14716 10848 14720
rect 10784 14660 10788 14716
rect 10788 14660 10844 14716
rect 10844 14660 10848 14716
rect 10784 14656 10848 14660
rect 10864 14716 10928 14720
rect 10864 14660 10868 14716
rect 10868 14660 10924 14716
rect 10924 14660 10928 14716
rect 10864 14656 10928 14660
rect 10944 14716 11008 14720
rect 10944 14660 10948 14716
rect 10948 14660 11004 14716
rect 11004 14660 11008 14716
rect 10944 14656 11008 14660
rect 11024 14716 11088 14720
rect 11024 14660 11028 14716
rect 11028 14660 11084 14716
rect 11084 14660 11088 14716
rect 11024 14656 11088 14660
rect 14717 14716 14781 14720
rect 14717 14660 14721 14716
rect 14721 14660 14777 14716
rect 14777 14660 14781 14716
rect 14717 14656 14781 14660
rect 14797 14716 14861 14720
rect 14797 14660 14801 14716
rect 14801 14660 14857 14716
rect 14857 14660 14861 14716
rect 14797 14656 14861 14660
rect 14877 14716 14941 14720
rect 14877 14660 14881 14716
rect 14881 14660 14937 14716
rect 14937 14660 14941 14716
rect 14877 14656 14941 14660
rect 14957 14716 15021 14720
rect 14957 14660 14961 14716
rect 14961 14660 15017 14716
rect 15017 14660 15021 14716
rect 14957 14656 15021 14660
rect 4884 14172 4948 14176
rect 4884 14116 4888 14172
rect 4888 14116 4944 14172
rect 4944 14116 4948 14172
rect 4884 14112 4948 14116
rect 4964 14172 5028 14176
rect 4964 14116 4968 14172
rect 4968 14116 5024 14172
rect 5024 14116 5028 14172
rect 4964 14112 5028 14116
rect 5044 14172 5108 14176
rect 5044 14116 5048 14172
rect 5048 14116 5104 14172
rect 5104 14116 5108 14172
rect 5044 14112 5108 14116
rect 5124 14172 5188 14176
rect 5124 14116 5128 14172
rect 5128 14116 5184 14172
rect 5184 14116 5188 14172
rect 5124 14112 5188 14116
rect 8817 14172 8881 14176
rect 8817 14116 8821 14172
rect 8821 14116 8877 14172
rect 8877 14116 8881 14172
rect 8817 14112 8881 14116
rect 8897 14172 8961 14176
rect 8897 14116 8901 14172
rect 8901 14116 8957 14172
rect 8957 14116 8961 14172
rect 8897 14112 8961 14116
rect 8977 14172 9041 14176
rect 8977 14116 8981 14172
rect 8981 14116 9037 14172
rect 9037 14116 9041 14172
rect 8977 14112 9041 14116
rect 9057 14172 9121 14176
rect 9057 14116 9061 14172
rect 9061 14116 9117 14172
rect 9117 14116 9121 14172
rect 9057 14112 9121 14116
rect 12750 14172 12814 14176
rect 12750 14116 12754 14172
rect 12754 14116 12810 14172
rect 12810 14116 12814 14172
rect 12750 14112 12814 14116
rect 12830 14172 12894 14176
rect 12830 14116 12834 14172
rect 12834 14116 12890 14172
rect 12890 14116 12894 14172
rect 12830 14112 12894 14116
rect 12910 14172 12974 14176
rect 12910 14116 12914 14172
rect 12914 14116 12970 14172
rect 12970 14116 12974 14172
rect 12910 14112 12974 14116
rect 12990 14172 13054 14176
rect 12990 14116 12994 14172
rect 12994 14116 13050 14172
rect 13050 14116 13054 14172
rect 12990 14112 13054 14116
rect 16683 14172 16747 14176
rect 16683 14116 16687 14172
rect 16687 14116 16743 14172
rect 16743 14116 16747 14172
rect 16683 14112 16747 14116
rect 16763 14172 16827 14176
rect 16763 14116 16767 14172
rect 16767 14116 16823 14172
rect 16823 14116 16827 14172
rect 16763 14112 16827 14116
rect 16843 14172 16907 14176
rect 16843 14116 16847 14172
rect 16847 14116 16903 14172
rect 16903 14116 16907 14172
rect 16843 14112 16907 14116
rect 16923 14172 16987 14176
rect 16923 14116 16927 14172
rect 16927 14116 16983 14172
rect 16983 14116 16987 14172
rect 16923 14112 16987 14116
rect 2918 13628 2982 13632
rect 2918 13572 2922 13628
rect 2922 13572 2978 13628
rect 2978 13572 2982 13628
rect 2918 13568 2982 13572
rect 2998 13628 3062 13632
rect 2998 13572 3002 13628
rect 3002 13572 3058 13628
rect 3058 13572 3062 13628
rect 2998 13568 3062 13572
rect 3078 13628 3142 13632
rect 3078 13572 3082 13628
rect 3082 13572 3138 13628
rect 3138 13572 3142 13628
rect 3078 13568 3142 13572
rect 3158 13628 3222 13632
rect 3158 13572 3162 13628
rect 3162 13572 3218 13628
rect 3218 13572 3222 13628
rect 3158 13568 3222 13572
rect 6851 13628 6915 13632
rect 6851 13572 6855 13628
rect 6855 13572 6911 13628
rect 6911 13572 6915 13628
rect 6851 13568 6915 13572
rect 6931 13628 6995 13632
rect 6931 13572 6935 13628
rect 6935 13572 6991 13628
rect 6991 13572 6995 13628
rect 6931 13568 6995 13572
rect 7011 13628 7075 13632
rect 7011 13572 7015 13628
rect 7015 13572 7071 13628
rect 7071 13572 7075 13628
rect 7011 13568 7075 13572
rect 7091 13628 7155 13632
rect 7091 13572 7095 13628
rect 7095 13572 7151 13628
rect 7151 13572 7155 13628
rect 7091 13568 7155 13572
rect 10784 13628 10848 13632
rect 10784 13572 10788 13628
rect 10788 13572 10844 13628
rect 10844 13572 10848 13628
rect 10784 13568 10848 13572
rect 10864 13628 10928 13632
rect 10864 13572 10868 13628
rect 10868 13572 10924 13628
rect 10924 13572 10928 13628
rect 10864 13568 10928 13572
rect 10944 13628 11008 13632
rect 10944 13572 10948 13628
rect 10948 13572 11004 13628
rect 11004 13572 11008 13628
rect 10944 13568 11008 13572
rect 11024 13628 11088 13632
rect 11024 13572 11028 13628
rect 11028 13572 11084 13628
rect 11084 13572 11088 13628
rect 11024 13568 11088 13572
rect 14717 13628 14781 13632
rect 14717 13572 14721 13628
rect 14721 13572 14777 13628
rect 14777 13572 14781 13628
rect 14717 13568 14781 13572
rect 14797 13628 14861 13632
rect 14797 13572 14801 13628
rect 14801 13572 14857 13628
rect 14857 13572 14861 13628
rect 14797 13568 14861 13572
rect 14877 13628 14941 13632
rect 14877 13572 14881 13628
rect 14881 13572 14937 13628
rect 14937 13572 14941 13628
rect 14877 13568 14941 13572
rect 14957 13628 15021 13632
rect 14957 13572 14961 13628
rect 14961 13572 15017 13628
rect 15017 13572 15021 13628
rect 14957 13568 15021 13572
rect 4884 13084 4948 13088
rect 4884 13028 4888 13084
rect 4888 13028 4944 13084
rect 4944 13028 4948 13084
rect 4884 13024 4948 13028
rect 4964 13084 5028 13088
rect 4964 13028 4968 13084
rect 4968 13028 5024 13084
rect 5024 13028 5028 13084
rect 4964 13024 5028 13028
rect 5044 13084 5108 13088
rect 5044 13028 5048 13084
rect 5048 13028 5104 13084
rect 5104 13028 5108 13084
rect 5044 13024 5108 13028
rect 5124 13084 5188 13088
rect 5124 13028 5128 13084
rect 5128 13028 5184 13084
rect 5184 13028 5188 13084
rect 5124 13024 5188 13028
rect 8817 13084 8881 13088
rect 8817 13028 8821 13084
rect 8821 13028 8877 13084
rect 8877 13028 8881 13084
rect 8817 13024 8881 13028
rect 8897 13084 8961 13088
rect 8897 13028 8901 13084
rect 8901 13028 8957 13084
rect 8957 13028 8961 13084
rect 8897 13024 8961 13028
rect 8977 13084 9041 13088
rect 8977 13028 8981 13084
rect 8981 13028 9037 13084
rect 9037 13028 9041 13084
rect 8977 13024 9041 13028
rect 9057 13084 9121 13088
rect 9057 13028 9061 13084
rect 9061 13028 9117 13084
rect 9117 13028 9121 13084
rect 9057 13024 9121 13028
rect 12750 13084 12814 13088
rect 12750 13028 12754 13084
rect 12754 13028 12810 13084
rect 12810 13028 12814 13084
rect 12750 13024 12814 13028
rect 12830 13084 12894 13088
rect 12830 13028 12834 13084
rect 12834 13028 12890 13084
rect 12890 13028 12894 13084
rect 12830 13024 12894 13028
rect 12910 13084 12974 13088
rect 12910 13028 12914 13084
rect 12914 13028 12970 13084
rect 12970 13028 12974 13084
rect 12910 13024 12974 13028
rect 12990 13084 13054 13088
rect 12990 13028 12994 13084
rect 12994 13028 13050 13084
rect 13050 13028 13054 13084
rect 12990 13024 13054 13028
rect 16683 13084 16747 13088
rect 16683 13028 16687 13084
rect 16687 13028 16743 13084
rect 16743 13028 16747 13084
rect 16683 13024 16747 13028
rect 16763 13084 16827 13088
rect 16763 13028 16767 13084
rect 16767 13028 16823 13084
rect 16823 13028 16827 13084
rect 16763 13024 16827 13028
rect 16843 13084 16907 13088
rect 16843 13028 16847 13084
rect 16847 13028 16903 13084
rect 16903 13028 16907 13084
rect 16843 13024 16907 13028
rect 16923 13084 16987 13088
rect 16923 13028 16927 13084
rect 16927 13028 16983 13084
rect 16983 13028 16987 13084
rect 16923 13024 16987 13028
rect 2918 12540 2982 12544
rect 2918 12484 2922 12540
rect 2922 12484 2978 12540
rect 2978 12484 2982 12540
rect 2918 12480 2982 12484
rect 2998 12540 3062 12544
rect 2998 12484 3002 12540
rect 3002 12484 3058 12540
rect 3058 12484 3062 12540
rect 2998 12480 3062 12484
rect 3078 12540 3142 12544
rect 3078 12484 3082 12540
rect 3082 12484 3138 12540
rect 3138 12484 3142 12540
rect 3078 12480 3142 12484
rect 3158 12540 3222 12544
rect 3158 12484 3162 12540
rect 3162 12484 3218 12540
rect 3218 12484 3222 12540
rect 3158 12480 3222 12484
rect 6851 12540 6915 12544
rect 6851 12484 6855 12540
rect 6855 12484 6911 12540
rect 6911 12484 6915 12540
rect 6851 12480 6915 12484
rect 6931 12540 6995 12544
rect 6931 12484 6935 12540
rect 6935 12484 6991 12540
rect 6991 12484 6995 12540
rect 6931 12480 6995 12484
rect 7011 12540 7075 12544
rect 7011 12484 7015 12540
rect 7015 12484 7071 12540
rect 7071 12484 7075 12540
rect 7011 12480 7075 12484
rect 7091 12540 7155 12544
rect 7091 12484 7095 12540
rect 7095 12484 7151 12540
rect 7151 12484 7155 12540
rect 7091 12480 7155 12484
rect 10784 12540 10848 12544
rect 10784 12484 10788 12540
rect 10788 12484 10844 12540
rect 10844 12484 10848 12540
rect 10784 12480 10848 12484
rect 10864 12540 10928 12544
rect 10864 12484 10868 12540
rect 10868 12484 10924 12540
rect 10924 12484 10928 12540
rect 10864 12480 10928 12484
rect 10944 12540 11008 12544
rect 10944 12484 10948 12540
rect 10948 12484 11004 12540
rect 11004 12484 11008 12540
rect 10944 12480 11008 12484
rect 11024 12540 11088 12544
rect 11024 12484 11028 12540
rect 11028 12484 11084 12540
rect 11084 12484 11088 12540
rect 11024 12480 11088 12484
rect 14717 12540 14781 12544
rect 14717 12484 14721 12540
rect 14721 12484 14777 12540
rect 14777 12484 14781 12540
rect 14717 12480 14781 12484
rect 14797 12540 14861 12544
rect 14797 12484 14801 12540
rect 14801 12484 14857 12540
rect 14857 12484 14861 12540
rect 14797 12480 14861 12484
rect 14877 12540 14941 12544
rect 14877 12484 14881 12540
rect 14881 12484 14937 12540
rect 14937 12484 14941 12540
rect 14877 12480 14941 12484
rect 14957 12540 15021 12544
rect 14957 12484 14961 12540
rect 14961 12484 15017 12540
rect 15017 12484 15021 12540
rect 14957 12480 15021 12484
rect 4884 11996 4948 12000
rect 4884 11940 4888 11996
rect 4888 11940 4944 11996
rect 4944 11940 4948 11996
rect 4884 11936 4948 11940
rect 4964 11996 5028 12000
rect 4964 11940 4968 11996
rect 4968 11940 5024 11996
rect 5024 11940 5028 11996
rect 4964 11936 5028 11940
rect 5044 11996 5108 12000
rect 5044 11940 5048 11996
rect 5048 11940 5104 11996
rect 5104 11940 5108 11996
rect 5044 11936 5108 11940
rect 5124 11996 5188 12000
rect 5124 11940 5128 11996
rect 5128 11940 5184 11996
rect 5184 11940 5188 11996
rect 5124 11936 5188 11940
rect 8817 11996 8881 12000
rect 8817 11940 8821 11996
rect 8821 11940 8877 11996
rect 8877 11940 8881 11996
rect 8817 11936 8881 11940
rect 8897 11996 8961 12000
rect 8897 11940 8901 11996
rect 8901 11940 8957 11996
rect 8957 11940 8961 11996
rect 8897 11936 8961 11940
rect 8977 11996 9041 12000
rect 8977 11940 8981 11996
rect 8981 11940 9037 11996
rect 9037 11940 9041 11996
rect 8977 11936 9041 11940
rect 9057 11996 9121 12000
rect 9057 11940 9061 11996
rect 9061 11940 9117 11996
rect 9117 11940 9121 11996
rect 9057 11936 9121 11940
rect 12750 11996 12814 12000
rect 12750 11940 12754 11996
rect 12754 11940 12810 11996
rect 12810 11940 12814 11996
rect 12750 11936 12814 11940
rect 12830 11996 12894 12000
rect 12830 11940 12834 11996
rect 12834 11940 12890 11996
rect 12890 11940 12894 11996
rect 12830 11936 12894 11940
rect 12910 11996 12974 12000
rect 12910 11940 12914 11996
rect 12914 11940 12970 11996
rect 12970 11940 12974 11996
rect 12910 11936 12974 11940
rect 12990 11996 13054 12000
rect 12990 11940 12994 11996
rect 12994 11940 13050 11996
rect 13050 11940 13054 11996
rect 12990 11936 13054 11940
rect 16683 11996 16747 12000
rect 16683 11940 16687 11996
rect 16687 11940 16743 11996
rect 16743 11940 16747 11996
rect 16683 11936 16747 11940
rect 16763 11996 16827 12000
rect 16763 11940 16767 11996
rect 16767 11940 16823 11996
rect 16823 11940 16827 11996
rect 16763 11936 16827 11940
rect 16843 11996 16907 12000
rect 16843 11940 16847 11996
rect 16847 11940 16903 11996
rect 16903 11940 16907 11996
rect 16843 11936 16907 11940
rect 16923 11996 16987 12000
rect 16923 11940 16927 11996
rect 16927 11940 16983 11996
rect 16983 11940 16987 11996
rect 16923 11936 16987 11940
rect 2918 11452 2982 11456
rect 2918 11396 2922 11452
rect 2922 11396 2978 11452
rect 2978 11396 2982 11452
rect 2918 11392 2982 11396
rect 2998 11452 3062 11456
rect 2998 11396 3002 11452
rect 3002 11396 3058 11452
rect 3058 11396 3062 11452
rect 2998 11392 3062 11396
rect 3078 11452 3142 11456
rect 3078 11396 3082 11452
rect 3082 11396 3138 11452
rect 3138 11396 3142 11452
rect 3078 11392 3142 11396
rect 3158 11452 3222 11456
rect 3158 11396 3162 11452
rect 3162 11396 3218 11452
rect 3218 11396 3222 11452
rect 3158 11392 3222 11396
rect 6851 11452 6915 11456
rect 6851 11396 6855 11452
rect 6855 11396 6911 11452
rect 6911 11396 6915 11452
rect 6851 11392 6915 11396
rect 6931 11452 6995 11456
rect 6931 11396 6935 11452
rect 6935 11396 6991 11452
rect 6991 11396 6995 11452
rect 6931 11392 6995 11396
rect 7011 11452 7075 11456
rect 7011 11396 7015 11452
rect 7015 11396 7071 11452
rect 7071 11396 7075 11452
rect 7011 11392 7075 11396
rect 7091 11452 7155 11456
rect 7091 11396 7095 11452
rect 7095 11396 7151 11452
rect 7151 11396 7155 11452
rect 7091 11392 7155 11396
rect 10784 11452 10848 11456
rect 10784 11396 10788 11452
rect 10788 11396 10844 11452
rect 10844 11396 10848 11452
rect 10784 11392 10848 11396
rect 10864 11452 10928 11456
rect 10864 11396 10868 11452
rect 10868 11396 10924 11452
rect 10924 11396 10928 11452
rect 10864 11392 10928 11396
rect 10944 11452 11008 11456
rect 10944 11396 10948 11452
rect 10948 11396 11004 11452
rect 11004 11396 11008 11452
rect 10944 11392 11008 11396
rect 11024 11452 11088 11456
rect 11024 11396 11028 11452
rect 11028 11396 11084 11452
rect 11084 11396 11088 11452
rect 11024 11392 11088 11396
rect 14717 11452 14781 11456
rect 14717 11396 14721 11452
rect 14721 11396 14777 11452
rect 14777 11396 14781 11452
rect 14717 11392 14781 11396
rect 14797 11452 14861 11456
rect 14797 11396 14801 11452
rect 14801 11396 14857 11452
rect 14857 11396 14861 11452
rect 14797 11392 14861 11396
rect 14877 11452 14941 11456
rect 14877 11396 14881 11452
rect 14881 11396 14937 11452
rect 14937 11396 14941 11452
rect 14877 11392 14941 11396
rect 14957 11452 15021 11456
rect 14957 11396 14961 11452
rect 14961 11396 15017 11452
rect 15017 11396 15021 11452
rect 14957 11392 15021 11396
rect 4884 10908 4948 10912
rect 4884 10852 4888 10908
rect 4888 10852 4944 10908
rect 4944 10852 4948 10908
rect 4884 10848 4948 10852
rect 4964 10908 5028 10912
rect 4964 10852 4968 10908
rect 4968 10852 5024 10908
rect 5024 10852 5028 10908
rect 4964 10848 5028 10852
rect 5044 10908 5108 10912
rect 5044 10852 5048 10908
rect 5048 10852 5104 10908
rect 5104 10852 5108 10908
rect 5044 10848 5108 10852
rect 5124 10908 5188 10912
rect 5124 10852 5128 10908
rect 5128 10852 5184 10908
rect 5184 10852 5188 10908
rect 5124 10848 5188 10852
rect 8817 10908 8881 10912
rect 8817 10852 8821 10908
rect 8821 10852 8877 10908
rect 8877 10852 8881 10908
rect 8817 10848 8881 10852
rect 8897 10908 8961 10912
rect 8897 10852 8901 10908
rect 8901 10852 8957 10908
rect 8957 10852 8961 10908
rect 8897 10848 8961 10852
rect 8977 10908 9041 10912
rect 8977 10852 8981 10908
rect 8981 10852 9037 10908
rect 9037 10852 9041 10908
rect 8977 10848 9041 10852
rect 9057 10908 9121 10912
rect 9057 10852 9061 10908
rect 9061 10852 9117 10908
rect 9117 10852 9121 10908
rect 9057 10848 9121 10852
rect 12750 10908 12814 10912
rect 12750 10852 12754 10908
rect 12754 10852 12810 10908
rect 12810 10852 12814 10908
rect 12750 10848 12814 10852
rect 12830 10908 12894 10912
rect 12830 10852 12834 10908
rect 12834 10852 12890 10908
rect 12890 10852 12894 10908
rect 12830 10848 12894 10852
rect 12910 10908 12974 10912
rect 12910 10852 12914 10908
rect 12914 10852 12970 10908
rect 12970 10852 12974 10908
rect 12910 10848 12974 10852
rect 12990 10908 13054 10912
rect 12990 10852 12994 10908
rect 12994 10852 13050 10908
rect 13050 10852 13054 10908
rect 12990 10848 13054 10852
rect 16683 10908 16747 10912
rect 16683 10852 16687 10908
rect 16687 10852 16743 10908
rect 16743 10852 16747 10908
rect 16683 10848 16747 10852
rect 16763 10908 16827 10912
rect 16763 10852 16767 10908
rect 16767 10852 16823 10908
rect 16823 10852 16827 10908
rect 16763 10848 16827 10852
rect 16843 10908 16907 10912
rect 16843 10852 16847 10908
rect 16847 10852 16903 10908
rect 16903 10852 16907 10908
rect 16843 10848 16907 10852
rect 16923 10908 16987 10912
rect 16923 10852 16927 10908
rect 16927 10852 16983 10908
rect 16983 10852 16987 10908
rect 16923 10848 16987 10852
rect 2918 10364 2982 10368
rect 2918 10308 2922 10364
rect 2922 10308 2978 10364
rect 2978 10308 2982 10364
rect 2918 10304 2982 10308
rect 2998 10364 3062 10368
rect 2998 10308 3002 10364
rect 3002 10308 3058 10364
rect 3058 10308 3062 10364
rect 2998 10304 3062 10308
rect 3078 10364 3142 10368
rect 3078 10308 3082 10364
rect 3082 10308 3138 10364
rect 3138 10308 3142 10364
rect 3078 10304 3142 10308
rect 3158 10364 3222 10368
rect 3158 10308 3162 10364
rect 3162 10308 3218 10364
rect 3218 10308 3222 10364
rect 3158 10304 3222 10308
rect 6851 10364 6915 10368
rect 6851 10308 6855 10364
rect 6855 10308 6911 10364
rect 6911 10308 6915 10364
rect 6851 10304 6915 10308
rect 6931 10364 6995 10368
rect 6931 10308 6935 10364
rect 6935 10308 6991 10364
rect 6991 10308 6995 10364
rect 6931 10304 6995 10308
rect 7011 10364 7075 10368
rect 7011 10308 7015 10364
rect 7015 10308 7071 10364
rect 7071 10308 7075 10364
rect 7011 10304 7075 10308
rect 7091 10364 7155 10368
rect 7091 10308 7095 10364
rect 7095 10308 7151 10364
rect 7151 10308 7155 10364
rect 7091 10304 7155 10308
rect 10784 10364 10848 10368
rect 10784 10308 10788 10364
rect 10788 10308 10844 10364
rect 10844 10308 10848 10364
rect 10784 10304 10848 10308
rect 10864 10364 10928 10368
rect 10864 10308 10868 10364
rect 10868 10308 10924 10364
rect 10924 10308 10928 10364
rect 10864 10304 10928 10308
rect 10944 10364 11008 10368
rect 10944 10308 10948 10364
rect 10948 10308 11004 10364
rect 11004 10308 11008 10364
rect 10944 10304 11008 10308
rect 11024 10364 11088 10368
rect 11024 10308 11028 10364
rect 11028 10308 11084 10364
rect 11084 10308 11088 10364
rect 11024 10304 11088 10308
rect 14717 10364 14781 10368
rect 14717 10308 14721 10364
rect 14721 10308 14777 10364
rect 14777 10308 14781 10364
rect 14717 10304 14781 10308
rect 14797 10364 14861 10368
rect 14797 10308 14801 10364
rect 14801 10308 14857 10364
rect 14857 10308 14861 10364
rect 14797 10304 14861 10308
rect 14877 10364 14941 10368
rect 14877 10308 14881 10364
rect 14881 10308 14937 10364
rect 14937 10308 14941 10364
rect 14877 10304 14941 10308
rect 14957 10364 15021 10368
rect 14957 10308 14961 10364
rect 14961 10308 15017 10364
rect 15017 10308 15021 10364
rect 14957 10304 15021 10308
rect 4884 9820 4948 9824
rect 4884 9764 4888 9820
rect 4888 9764 4944 9820
rect 4944 9764 4948 9820
rect 4884 9760 4948 9764
rect 4964 9820 5028 9824
rect 4964 9764 4968 9820
rect 4968 9764 5024 9820
rect 5024 9764 5028 9820
rect 4964 9760 5028 9764
rect 5044 9820 5108 9824
rect 5044 9764 5048 9820
rect 5048 9764 5104 9820
rect 5104 9764 5108 9820
rect 5044 9760 5108 9764
rect 5124 9820 5188 9824
rect 5124 9764 5128 9820
rect 5128 9764 5184 9820
rect 5184 9764 5188 9820
rect 5124 9760 5188 9764
rect 8817 9820 8881 9824
rect 8817 9764 8821 9820
rect 8821 9764 8877 9820
rect 8877 9764 8881 9820
rect 8817 9760 8881 9764
rect 8897 9820 8961 9824
rect 8897 9764 8901 9820
rect 8901 9764 8957 9820
rect 8957 9764 8961 9820
rect 8897 9760 8961 9764
rect 8977 9820 9041 9824
rect 8977 9764 8981 9820
rect 8981 9764 9037 9820
rect 9037 9764 9041 9820
rect 8977 9760 9041 9764
rect 9057 9820 9121 9824
rect 9057 9764 9061 9820
rect 9061 9764 9117 9820
rect 9117 9764 9121 9820
rect 9057 9760 9121 9764
rect 12750 9820 12814 9824
rect 12750 9764 12754 9820
rect 12754 9764 12810 9820
rect 12810 9764 12814 9820
rect 12750 9760 12814 9764
rect 12830 9820 12894 9824
rect 12830 9764 12834 9820
rect 12834 9764 12890 9820
rect 12890 9764 12894 9820
rect 12830 9760 12894 9764
rect 12910 9820 12974 9824
rect 12910 9764 12914 9820
rect 12914 9764 12970 9820
rect 12970 9764 12974 9820
rect 12910 9760 12974 9764
rect 12990 9820 13054 9824
rect 12990 9764 12994 9820
rect 12994 9764 13050 9820
rect 13050 9764 13054 9820
rect 12990 9760 13054 9764
rect 16683 9820 16747 9824
rect 16683 9764 16687 9820
rect 16687 9764 16743 9820
rect 16743 9764 16747 9820
rect 16683 9760 16747 9764
rect 16763 9820 16827 9824
rect 16763 9764 16767 9820
rect 16767 9764 16823 9820
rect 16823 9764 16827 9820
rect 16763 9760 16827 9764
rect 16843 9820 16907 9824
rect 16843 9764 16847 9820
rect 16847 9764 16903 9820
rect 16903 9764 16907 9820
rect 16843 9760 16907 9764
rect 16923 9820 16987 9824
rect 16923 9764 16927 9820
rect 16927 9764 16983 9820
rect 16983 9764 16987 9820
rect 16923 9760 16987 9764
rect 2918 9276 2982 9280
rect 2918 9220 2922 9276
rect 2922 9220 2978 9276
rect 2978 9220 2982 9276
rect 2918 9216 2982 9220
rect 2998 9276 3062 9280
rect 2998 9220 3002 9276
rect 3002 9220 3058 9276
rect 3058 9220 3062 9276
rect 2998 9216 3062 9220
rect 3078 9276 3142 9280
rect 3078 9220 3082 9276
rect 3082 9220 3138 9276
rect 3138 9220 3142 9276
rect 3078 9216 3142 9220
rect 3158 9276 3222 9280
rect 3158 9220 3162 9276
rect 3162 9220 3218 9276
rect 3218 9220 3222 9276
rect 3158 9216 3222 9220
rect 6851 9276 6915 9280
rect 6851 9220 6855 9276
rect 6855 9220 6911 9276
rect 6911 9220 6915 9276
rect 6851 9216 6915 9220
rect 6931 9276 6995 9280
rect 6931 9220 6935 9276
rect 6935 9220 6991 9276
rect 6991 9220 6995 9276
rect 6931 9216 6995 9220
rect 7011 9276 7075 9280
rect 7011 9220 7015 9276
rect 7015 9220 7071 9276
rect 7071 9220 7075 9276
rect 7011 9216 7075 9220
rect 7091 9276 7155 9280
rect 7091 9220 7095 9276
rect 7095 9220 7151 9276
rect 7151 9220 7155 9276
rect 7091 9216 7155 9220
rect 10784 9276 10848 9280
rect 10784 9220 10788 9276
rect 10788 9220 10844 9276
rect 10844 9220 10848 9276
rect 10784 9216 10848 9220
rect 10864 9276 10928 9280
rect 10864 9220 10868 9276
rect 10868 9220 10924 9276
rect 10924 9220 10928 9276
rect 10864 9216 10928 9220
rect 10944 9276 11008 9280
rect 10944 9220 10948 9276
rect 10948 9220 11004 9276
rect 11004 9220 11008 9276
rect 10944 9216 11008 9220
rect 11024 9276 11088 9280
rect 11024 9220 11028 9276
rect 11028 9220 11084 9276
rect 11084 9220 11088 9276
rect 11024 9216 11088 9220
rect 14717 9276 14781 9280
rect 14717 9220 14721 9276
rect 14721 9220 14777 9276
rect 14777 9220 14781 9276
rect 14717 9216 14781 9220
rect 14797 9276 14861 9280
rect 14797 9220 14801 9276
rect 14801 9220 14857 9276
rect 14857 9220 14861 9276
rect 14797 9216 14861 9220
rect 14877 9276 14941 9280
rect 14877 9220 14881 9276
rect 14881 9220 14937 9276
rect 14937 9220 14941 9276
rect 14877 9216 14941 9220
rect 14957 9276 15021 9280
rect 14957 9220 14961 9276
rect 14961 9220 15017 9276
rect 15017 9220 15021 9276
rect 14957 9216 15021 9220
rect 4884 8732 4948 8736
rect 4884 8676 4888 8732
rect 4888 8676 4944 8732
rect 4944 8676 4948 8732
rect 4884 8672 4948 8676
rect 4964 8732 5028 8736
rect 4964 8676 4968 8732
rect 4968 8676 5024 8732
rect 5024 8676 5028 8732
rect 4964 8672 5028 8676
rect 5044 8732 5108 8736
rect 5044 8676 5048 8732
rect 5048 8676 5104 8732
rect 5104 8676 5108 8732
rect 5044 8672 5108 8676
rect 5124 8732 5188 8736
rect 5124 8676 5128 8732
rect 5128 8676 5184 8732
rect 5184 8676 5188 8732
rect 5124 8672 5188 8676
rect 8817 8732 8881 8736
rect 8817 8676 8821 8732
rect 8821 8676 8877 8732
rect 8877 8676 8881 8732
rect 8817 8672 8881 8676
rect 8897 8732 8961 8736
rect 8897 8676 8901 8732
rect 8901 8676 8957 8732
rect 8957 8676 8961 8732
rect 8897 8672 8961 8676
rect 8977 8732 9041 8736
rect 8977 8676 8981 8732
rect 8981 8676 9037 8732
rect 9037 8676 9041 8732
rect 8977 8672 9041 8676
rect 9057 8732 9121 8736
rect 9057 8676 9061 8732
rect 9061 8676 9117 8732
rect 9117 8676 9121 8732
rect 9057 8672 9121 8676
rect 12750 8732 12814 8736
rect 12750 8676 12754 8732
rect 12754 8676 12810 8732
rect 12810 8676 12814 8732
rect 12750 8672 12814 8676
rect 12830 8732 12894 8736
rect 12830 8676 12834 8732
rect 12834 8676 12890 8732
rect 12890 8676 12894 8732
rect 12830 8672 12894 8676
rect 12910 8732 12974 8736
rect 12910 8676 12914 8732
rect 12914 8676 12970 8732
rect 12970 8676 12974 8732
rect 12910 8672 12974 8676
rect 12990 8732 13054 8736
rect 12990 8676 12994 8732
rect 12994 8676 13050 8732
rect 13050 8676 13054 8732
rect 12990 8672 13054 8676
rect 16683 8732 16747 8736
rect 16683 8676 16687 8732
rect 16687 8676 16743 8732
rect 16743 8676 16747 8732
rect 16683 8672 16747 8676
rect 16763 8732 16827 8736
rect 16763 8676 16767 8732
rect 16767 8676 16823 8732
rect 16823 8676 16827 8732
rect 16763 8672 16827 8676
rect 16843 8732 16907 8736
rect 16843 8676 16847 8732
rect 16847 8676 16903 8732
rect 16903 8676 16907 8732
rect 16843 8672 16907 8676
rect 16923 8732 16987 8736
rect 16923 8676 16927 8732
rect 16927 8676 16983 8732
rect 16983 8676 16987 8732
rect 16923 8672 16987 8676
rect 2918 8188 2982 8192
rect 2918 8132 2922 8188
rect 2922 8132 2978 8188
rect 2978 8132 2982 8188
rect 2918 8128 2982 8132
rect 2998 8188 3062 8192
rect 2998 8132 3002 8188
rect 3002 8132 3058 8188
rect 3058 8132 3062 8188
rect 2998 8128 3062 8132
rect 3078 8188 3142 8192
rect 3078 8132 3082 8188
rect 3082 8132 3138 8188
rect 3138 8132 3142 8188
rect 3078 8128 3142 8132
rect 3158 8188 3222 8192
rect 3158 8132 3162 8188
rect 3162 8132 3218 8188
rect 3218 8132 3222 8188
rect 3158 8128 3222 8132
rect 6851 8188 6915 8192
rect 6851 8132 6855 8188
rect 6855 8132 6911 8188
rect 6911 8132 6915 8188
rect 6851 8128 6915 8132
rect 6931 8188 6995 8192
rect 6931 8132 6935 8188
rect 6935 8132 6991 8188
rect 6991 8132 6995 8188
rect 6931 8128 6995 8132
rect 7011 8188 7075 8192
rect 7011 8132 7015 8188
rect 7015 8132 7071 8188
rect 7071 8132 7075 8188
rect 7011 8128 7075 8132
rect 7091 8188 7155 8192
rect 7091 8132 7095 8188
rect 7095 8132 7151 8188
rect 7151 8132 7155 8188
rect 7091 8128 7155 8132
rect 10784 8188 10848 8192
rect 10784 8132 10788 8188
rect 10788 8132 10844 8188
rect 10844 8132 10848 8188
rect 10784 8128 10848 8132
rect 10864 8188 10928 8192
rect 10864 8132 10868 8188
rect 10868 8132 10924 8188
rect 10924 8132 10928 8188
rect 10864 8128 10928 8132
rect 10944 8188 11008 8192
rect 10944 8132 10948 8188
rect 10948 8132 11004 8188
rect 11004 8132 11008 8188
rect 10944 8128 11008 8132
rect 11024 8188 11088 8192
rect 11024 8132 11028 8188
rect 11028 8132 11084 8188
rect 11084 8132 11088 8188
rect 11024 8128 11088 8132
rect 14717 8188 14781 8192
rect 14717 8132 14721 8188
rect 14721 8132 14777 8188
rect 14777 8132 14781 8188
rect 14717 8128 14781 8132
rect 14797 8188 14861 8192
rect 14797 8132 14801 8188
rect 14801 8132 14857 8188
rect 14857 8132 14861 8188
rect 14797 8128 14861 8132
rect 14877 8188 14941 8192
rect 14877 8132 14881 8188
rect 14881 8132 14937 8188
rect 14937 8132 14941 8188
rect 14877 8128 14941 8132
rect 14957 8188 15021 8192
rect 14957 8132 14961 8188
rect 14961 8132 15017 8188
rect 15017 8132 15021 8188
rect 14957 8128 15021 8132
rect 4884 7644 4948 7648
rect 4884 7588 4888 7644
rect 4888 7588 4944 7644
rect 4944 7588 4948 7644
rect 4884 7584 4948 7588
rect 4964 7644 5028 7648
rect 4964 7588 4968 7644
rect 4968 7588 5024 7644
rect 5024 7588 5028 7644
rect 4964 7584 5028 7588
rect 5044 7644 5108 7648
rect 5044 7588 5048 7644
rect 5048 7588 5104 7644
rect 5104 7588 5108 7644
rect 5044 7584 5108 7588
rect 5124 7644 5188 7648
rect 5124 7588 5128 7644
rect 5128 7588 5184 7644
rect 5184 7588 5188 7644
rect 5124 7584 5188 7588
rect 8817 7644 8881 7648
rect 8817 7588 8821 7644
rect 8821 7588 8877 7644
rect 8877 7588 8881 7644
rect 8817 7584 8881 7588
rect 8897 7644 8961 7648
rect 8897 7588 8901 7644
rect 8901 7588 8957 7644
rect 8957 7588 8961 7644
rect 8897 7584 8961 7588
rect 8977 7644 9041 7648
rect 8977 7588 8981 7644
rect 8981 7588 9037 7644
rect 9037 7588 9041 7644
rect 8977 7584 9041 7588
rect 9057 7644 9121 7648
rect 9057 7588 9061 7644
rect 9061 7588 9117 7644
rect 9117 7588 9121 7644
rect 9057 7584 9121 7588
rect 12750 7644 12814 7648
rect 12750 7588 12754 7644
rect 12754 7588 12810 7644
rect 12810 7588 12814 7644
rect 12750 7584 12814 7588
rect 12830 7644 12894 7648
rect 12830 7588 12834 7644
rect 12834 7588 12890 7644
rect 12890 7588 12894 7644
rect 12830 7584 12894 7588
rect 12910 7644 12974 7648
rect 12910 7588 12914 7644
rect 12914 7588 12970 7644
rect 12970 7588 12974 7644
rect 12910 7584 12974 7588
rect 12990 7644 13054 7648
rect 12990 7588 12994 7644
rect 12994 7588 13050 7644
rect 13050 7588 13054 7644
rect 12990 7584 13054 7588
rect 16683 7644 16747 7648
rect 16683 7588 16687 7644
rect 16687 7588 16743 7644
rect 16743 7588 16747 7644
rect 16683 7584 16747 7588
rect 16763 7644 16827 7648
rect 16763 7588 16767 7644
rect 16767 7588 16823 7644
rect 16823 7588 16827 7644
rect 16763 7584 16827 7588
rect 16843 7644 16907 7648
rect 16843 7588 16847 7644
rect 16847 7588 16903 7644
rect 16903 7588 16907 7644
rect 16843 7584 16907 7588
rect 16923 7644 16987 7648
rect 16923 7588 16927 7644
rect 16927 7588 16983 7644
rect 16983 7588 16987 7644
rect 16923 7584 16987 7588
rect 2918 7100 2982 7104
rect 2918 7044 2922 7100
rect 2922 7044 2978 7100
rect 2978 7044 2982 7100
rect 2918 7040 2982 7044
rect 2998 7100 3062 7104
rect 2998 7044 3002 7100
rect 3002 7044 3058 7100
rect 3058 7044 3062 7100
rect 2998 7040 3062 7044
rect 3078 7100 3142 7104
rect 3078 7044 3082 7100
rect 3082 7044 3138 7100
rect 3138 7044 3142 7100
rect 3078 7040 3142 7044
rect 3158 7100 3222 7104
rect 3158 7044 3162 7100
rect 3162 7044 3218 7100
rect 3218 7044 3222 7100
rect 3158 7040 3222 7044
rect 6851 7100 6915 7104
rect 6851 7044 6855 7100
rect 6855 7044 6911 7100
rect 6911 7044 6915 7100
rect 6851 7040 6915 7044
rect 6931 7100 6995 7104
rect 6931 7044 6935 7100
rect 6935 7044 6991 7100
rect 6991 7044 6995 7100
rect 6931 7040 6995 7044
rect 7011 7100 7075 7104
rect 7011 7044 7015 7100
rect 7015 7044 7071 7100
rect 7071 7044 7075 7100
rect 7011 7040 7075 7044
rect 7091 7100 7155 7104
rect 7091 7044 7095 7100
rect 7095 7044 7151 7100
rect 7151 7044 7155 7100
rect 7091 7040 7155 7044
rect 10784 7100 10848 7104
rect 10784 7044 10788 7100
rect 10788 7044 10844 7100
rect 10844 7044 10848 7100
rect 10784 7040 10848 7044
rect 10864 7100 10928 7104
rect 10864 7044 10868 7100
rect 10868 7044 10924 7100
rect 10924 7044 10928 7100
rect 10864 7040 10928 7044
rect 10944 7100 11008 7104
rect 10944 7044 10948 7100
rect 10948 7044 11004 7100
rect 11004 7044 11008 7100
rect 10944 7040 11008 7044
rect 11024 7100 11088 7104
rect 11024 7044 11028 7100
rect 11028 7044 11084 7100
rect 11084 7044 11088 7100
rect 11024 7040 11088 7044
rect 14717 7100 14781 7104
rect 14717 7044 14721 7100
rect 14721 7044 14777 7100
rect 14777 7044 14781 7100
rect 14717 7040 14781 7044
rect 14797 7100 14861 7104
rect 14797 7044 14801 7100
rect 14801 7044 14857 7100
rect 14857 7044 14861 7100
rect 14797 7040 14861 7044
rect 14877 7100 14941 7104
rect 14877 7044 14881 7100
rect 14881 7044 14937 7100
rect 14937 7044 14941 7100
rect 14877 7040 14941 7044
rect 14957 7100 15021 7104
rect 14957 7044 14961 7100
rect 14961 7044 15017 7100
rect 15017 7044 15021 7100
rect 14957 7040 15021 7044
rect 4884 6556 4948 6560
rect 4884 6500 4888 6556
rect 4888 6500 4944 6556
rect 4944 6500 4948 6556
rect 4884 6496 4948 6500
rect 4964 6556 5028 6560
rect 4964 6500 4968 6556
rect 4968 6500 5024 6556
rect 5024 6500 5028 6556
rect 4964 6496 5028 6500
rect 5044 6556 5108 6560
rect 5044 6500 5048 6556
rect 5048 6500 5104 6556
rect 5104 6500 5108 6556
rect 5044 6496 5108 6500
rect 5124 6556 5188 6560
rect 5124 6500 5128 6556
rect 5128 6500 5184 6556
rect 5184 6500 5188 6556
rect 5124 6496 5188 6500
rect 8817 6556 8881 6560
rect 8817 6500 8821 6556
rect 8821 6500 8877 6556
rect 8877 6500 8881 6556
rect 8817 6496 8881 6500
rect 8897 6556 8961 6560
rect 8897 6500 8901 6556
rect 8901 6500 8957 6556
rect 8957 6500 8961 6556
rect 8897 6496 8961 6500
rect 8977 6556 9041 6560
rect 8977 6500 8981 6556
rect 8981 6500 9037 6556
rect 9037 6500 9041 6556
rect 8977 6496 9041 6500
rect 9057 6556 9121 6560
rect 9057 6500 9061 6556
rect 9061 6500 9117 6556
rect 9117 6500 9121 6556
rect 9057 6496 9121 6500
rect 12750 6556 12814 6560
rect 12750 6500 12754 6556
rect 12754 6500 12810 6556
rect 12810 6500 12814 6556
rect 12750 6496 12814 6500
rect 12830 6556 12894 6560
rect 12830 6500 12834 6556
rect 12834 6500 12890 6556
rect 12890 6500 12894 6556
rect 12830 6496 12894 6500
rect 12910 6556 12974 6560
rect 12910 6500 12914 6556
rect 12914 6500 12970 6556
rect 12970 6500 12974 6556
rect 12910 6496 12974 6500
rect 12990 6556 13054 6560
rect 12990 6500 12994 6556
rect 12994 6500 13050 6556
rect 13050 6500 13054 6556
rect 12990 6496 13054 6500
rect 16683 6556 16747 6560
rect 16683 6500 16687 6556
rect 16687 6500 16743 6556
rect 16743 6500 16747 6556
rect 16683 6496 16747 6500
rect 16763 6556 16827 6560
rect 16763 6500 16767 6556
rect 16767 6500 16823 6556
rect 16823 6500 16827 6556
rect 16763 6496 16827 6500
rect 16843 6556 16907 6560
rect 16843 6500 16847 6556
rect 16847 6500 16903 6556
rect 16903 6500 16907 6556
rect 16843 6496 16907 6500
rect 16923 6556 16987 6560
rect 16923 6500 16927 6556
rect 16927 6500 16983 6556
rect 16983 6500 16987 6556
rect 16923 6496 16987 6500
rect 2918 6012 2982 6016
rect 2918 5956 2922 6012
rect 2922 5956 2978 6012
rect 2978 5956 2982 6012
rect 2918 5952 2982 5956
rect 2998 6012 3062 6016
rect 2998 5956 3002 6012
rect 3002 5956 3058 6012
rect 3058 5956 3062 6012
rect 2998 5952 3062 5956
rect 3078 6012 3142 6016
rect 3078 5956 3082 6012
rect 3082 5956 3138 6012
rect 3138 5956 3142 6012
rect 3078 5952 3142 5956
rect 3158 6012 3222 6016
rect 3158 5956 3162 6012
rect 3162 5956 3218 6012
rect 3218 5956 3222 6012
rect 3158 5952 3222 5956
rect 6851 6012 6915 6016
rect 6851 5956 6855 6012
rect 6855 5956 6911 6012
rect 6911 5956 6915 6012
rect 6851 5952 6915 5956
rect 6931 6012 6995 6016
rect 6931 5956 6935 6012
rect 6935 5956 6991 6012
rect 6991 5956 6995 6012
rect 6931 5952 6995 5956
rect 7011 6012 7075 6016
rect 7011 5956 7015 6012
rect 7015 5956 7071 6012
rect 7071 5956 7075 6012
rect 7011 5952 7075 5956
rect 7091 6012 7155 6016
rect 7091 5956 7095 6012
rect 7095 5956 7151 6012
rect 7151 5956 7155 6012
rect 7091 5952 7155 5956
rect 10784 6012 10848 6016
rect 10784 5956 10788 6012
rect 10788 5956 10844 6012
rect 10844 5956 10848 6012
rect 10784 5952 10848 5956
rect 10864 6012 10928 6016
rect 10864 5956 10868 6012
rect 10868 5956 10924 6012
rect 10924 5956 10928 6012
rect 10864 5952 10928 5956
rect 10944 6012 11008 6016
rect 10944 5956 10948 6012
rect 10948 5956 11004 6012
rect 11004 5956 11008 6012
rect 10944 5952 11008 5956
rect 11024 6012 11088 6016
rect 11024 5956 11028 6012
rect 11028 5956 11084 6012
rect 11084 5956 11088 6012
rect 11024 5952 11088 5956
rect 14717 6012 14781 6016
rect 14717 5956 14721 6012
rect 14721 5956 14777 6012
rect 14777 5956 14781 6012
rect 14717 5952 14781 5956
rect 14797 6012 14861 6016
rect 14797 5956 14801 6012
rect 14801 5956 14857 6012
rect 14857 5956 14861 6012
rect 14797 5952 14861 5956
rect 14877 6012 14941 6016
rect 14877 5956 14881 6012
rect 14881 5956 14937 6012
rect 14937 5956 14941 6012
rect 14877 5952 14941 5956
rect 14957 6012 15021 6016
rect 14957 5956 14961 6012
rect 14961 5956 15017 6012
rect 15017 5956 15021 6012
rect 14957 5952 15021 5956
rect 4884 5468 4948 5472
rect 4884 5412 4888 5468
rect 4888 5412 4944 5468
rect 4944 5412 4948 5468
rect 4884 5408 4948 5412
rect 4964 5468 5028 5472
rect 4964 5412 4968 5468
rect 4968 5412 5024 5468
rect 5024 5412 5028 5468
rect 4964 5408 5028 5412
rect 5044 5468 5108 5472
rect 5044 5412 5048 5468
rect 5048 5412 5104 5468
rect 5104 5412 5108 5468
rect 5044 5408 5108 5412
rect 5124 5468 5188 5472
rect 5124 5412 5128 5468
rect 5128 5412 5184 5468
rect 5184 5412 5188 5468
rect 5124 5408 5188 5412
rect 8817 5468 8881 5472
rect 8817 5412 8821 5468
rect 8821 5412 8877 5468
rect 8877 5412 8881 5468
rect 8817 5408 8881 5412
rect 8897 5468 8961 5472
rect 8897 5412 8901 5468
rect 8901 5412 8957 5468
rect 8957 5412 8961 5468
rect 8897 5408 8961 5412
rect 8977 5468 9041 5472
rect 8977 5412 8981 5468
rect 8981 5412 9037 5468
rect 9037 5412 9041 5468
rect 8977 5408 9041 5412
rect 9057 5468 9121 5472
rect 9057 5412 9061 5468
rect 9061 5412 9117 5468
rect 9117 5412 9121 5468
rect 9057 5408 9121 5412
rect 12750 5468 12814 5472
rect 12750 5412 12754 5468
rect 12754 5412 12810 5468
rect 12810 5412 12814 5468
rect 12750 5408 12814 5412
rect 12830 5468 12894 5472
rect 12830 5412 12834 5468
rect 12834 5412 12890 5468
rect 12890 5412 12894 5468
rect 12830 5408 12894 5412
rect 12910 5468 12974 5472
rect 12910 5412 12914 5468
rect 12914 5412 12970 5468
rect 12970 5412 12974 5468
rect 12910 5408 12974 5412
rect 12990 5468 13054 5472
rect 12990 5412 12994 5468
rect 12994 5412 13050 5468
rect 13050 5412 13054 5468
rect 12990 5408 13054 5412
rect 16683 5468 16747 5472
rect 16683 5412 16687 5468
rect 16687 5412 16743 5468
rect 16743 5412 16747 5468
rect 16683 5408 16747 5412
rect 16763 5468 16827 5472
rect 16763 5412 16767 5468
rect 16767 5412 16823 5468
rect 16823 5412 16827 5468
rect 16763 5408 16827 5412
rect 16843 5468 16907 5472
rect 16843 5412 16847 5468
rect 16847 5412 16903 5468
rect 16903 5412 16907 5468
rect 16843 5408 16907 5412
rect 16923 5468 16987 5472
rect 16923 5412 16927 5468
rect 16927 5412 16983 5468
rect 16983 5412 16987 5468
rect 16923 5408 16987 5412
rect 2918 4924 2982 4928
rect 2918 4868 2922 4924
rect 2922 4868 2978 4924
rect 2978 4868 2982 4924
rect 2918 4864 2982 4868
rect 2998 4924 3062 4928
rect 2998 4868 3002 4924
rect 3002 4868 3058 4924
rect 3058 4868 3062 4924
rect 2998 4864 3062 4868
rect 3078 4924 3142 4928
rect 3078 4868 3082 4924
rect 3082 4868 3138 4924
rect 3138 4868 3142 4924
rect 3078 4864 3142 4868
rect 3158 4924 3222 4928
rect 3158 4868 3162 4924
rect 3162 4868 3218 4924
rect 3218 4868 3222 4924
rect 3158 4864 3222 4868
rect 6851 4924 6915 4928
rect 6851 4868 6855 4924
rect 6855 4868 6911 4924
rect 6911 4868 6915 4924
rect 6851 4864 6915 4868
rect 6931 4924 6995 4928
rect 6931 4868 6935 4924
rect 6935 4868 6991 4924
rect 6991 4868 6995 4924
rect 6931 4864 6995 4868
rect 7011 4924 7075 4928
rect 7011 4868 7015 4924
rect 7015 4868 7071 4924
rect 7071 4868 7075 4924
rect 7011 4864 7075 4868
rect 7091 4924 7155 4928
rect 7091 4868 7095 4924
rect 7095 4868 7151 4924
rect 7151 4868 7155 4924
rect 7091 4864 7155 4868
rect 10784 4924 10848 4928
rect 10784 4868 10788 4924
rect 10788 4868 10844 4924
rect 10844 4868 10848 4924
rect 10784 4864 10848 4868
rect 10864 4924 10928 4928
rect 10864 4868 10868 4924
rect 10868 4868 10924 4924
rect 10924 4868 10928 4924
rect 10864 4864 10928 4868
rect 10944 4924 11008 4928
rect 10944 4868 10948 4924
rect 10948 4868 11004 4924
rect 11004 4868 11008 4924
rect 10944 4864 11008 4868
rect 11024 4924 11088 4928
rect 11024 4868 11028 4924
rect 11028 4868 11084 4924
rect 11084 4868 11088 4924
rect 11024 4864 11088 4868
rect 14717 4924 14781 4928
rect 14717 4868 14721 4924
rect 14721 4868 14777 4924
rect 14777 4868 14781 4924
rect 14717 4864 14781 4868
rect 14797 4924 14861 4928
rect 14797 4868 14801 4924
rect 14801 4868 14857 4924
rect 14857 4868 14861 4924
rect 14797 4864 14861 4868
rect 14877 4924 14941 4928
rect 14877 4868 14881 4924
rect 14881 4868 14937 4924
rect 14937 4868 14941 4924
rect 14877 4864 14941 4868
rect 14957 4924 15021 4928
rect 14957 4868 14961 4924
rect 14961 4868 15017 4924
rect 15017 4868 15021 4924
rect 14957 4864 15021 4868
rect 4884 4380 4948 4384
rect 4884 4324 4888 4380
rect 4888 4324 4944 4380
rect 4944 4324 4948 4380
rect 4884 4320 4948 4324
rect 4964 4380 5028 4384
rect 4964 4324 4968 4380
rect 4968 4324 5024 4380
rect 5024 4324 5028 4380
rect 4964 4320 5028 4324
rect 5044 4380 5108 4384
rect 5044 4324 5048 4380
rect 5048 4324 5104 4380
rect 5104 4324 5108 4380
rect 5044 4320 5108 4324
rect 5124 4380 5188 4384
rect 5124 4324 5128 4380
rect 5128 4324 5184 4380
rect 5184 4324 5188 4380
rect 5124 4320 5188 4324
rect 8817 4380 8881 4384
rect 8817 4324 8821 4380
rect 8821 4324 8877 4380
rect 8877 4324 8881 4380
rect 8817 4320 8881 4324
rect 8897 4380 8961 4384
rect 8897 4324 8901 4380
rect 8901 4324 8957 4380
rect 8957 4324 8961 4380
rect 8897 4320 8961 4324
rect 8977 4380 9041 4384
rect 8977 4324 8981 4380
rect 8981 4324 9037 4380
rect 9037 4324 9041 4380
rect 8977 4320 9041 4324
rect 9057 4380 9121 4384
rect 9057 4324 9061 4380
rect 9061 4324 9117 4380
rect 9117 4324 9121 4380
rect 9057 4320 9121 4324
rect 12750 4380 12814 4384
rect 12750 4324 12754 4380
rect 12754 4324 12810 4380
rect 12810 4324 12814 4380
rect 12750 4320 12814 4324
rect 12830 4380 12894 4384
rect 12830 4324 12834 4380
rect 12834 4324 12890 4380
rect 12890 4324 12894 4380
rect 12830 4320 12894 4324
rect 12910 4380 12974 4384
rect 12910 4324 12914 4380
rect 12914 4324 12970 4380
rect 12970 4324 12974 4380
rect 12910 4320 12974 4324
rect 12990 4380 13054 4384
rect 12990 4324 12994 4380
rect 12994 4324 13050 4380
rect 13050 4324 13054 4380
rect 12990 4320 13054 4324
rect 16683 4380 16747 4384
rect 16683 4324 16687 4380
rect 16687 4324 16743 4380
rect 16743 4324 16747 4380
rect 16683 4320 16747 4324
rect 16763 4380 16827 4384
rect 16763 4324 16767 4380
rect 16767 4324 16823 4380
rect 16823 4324 16827 4380
rect 16763 4320 16827 4324
rect 16843 4380 16907 4384
rect 16843 4324 16847 4380
rect 16847 4324 16903 4380
rect 16903 4324 16907 4380
rect 16843 4320 16907 4324
rect 16923 4380 16987 4384
rect 16923 4324 16927 4380
rect 16927 4324 16983 4380
rect 16983 4324 16987 4380
rect 16923 4320 16987 4324
rect 2918 3836 2982 3840
rect 2918 3780 2922 3836
rect 2922 3780 2978 3836
rect 2978 3780 2982 3836
rect 2918 3776 2982 3780
rect 2998 3836 3062 3840
rect 2998 3780 3002 3836
rect 3002 3780 3058 3836
rect 3058 3780 3062 3836
rect 2998 3776 3062 3780
rect 3078 3836 3142 3840
rect 3078 3780 3082 3836
rect 3082 3780 3138 3836
rect 3138 3780 3142 3836
rect 3078 3776 3142 3780
rect 3158 3836 3222 3840
rect 3158 3780 3162 3836
rect 3162 3780 3218 3836
rect 3218 3780 3222 3836
rect 3158 3776 3222 3780
rect 6851 3836 6915 3840
rect 6851 3780 6855 3836
rect 6855 3780 6911 3836
rect 6911 3780 6915 3836
rect 6851 3776 6915 3780
rect 6931 3836 6995 3840
rect 6931 3780 6935 3836
rect 6935 3780 6991 3836
rect 6991 3780 6995 3836
rect 6931 3776 6995 3780
rect 7011 3836 7075 3840
rect 7011 3780 7015 3836
rect 7015 3780 7071 3836
rect 7071 3780 7075 3836
rect 7011 3776 7075 3780
rect 7091 3836 7155 3840
rect 7091 3780 7095 3836
rect 7095 3780 7151 3836
rect 7151 3780 7155 3836
rect 7091 3776 7155 3780
rect 10784 3836 10848 3840
rect 10784 3780 10788 3836
rect 10788 3780 10844 3836
rect 10844 3780 10848 3836
rect 10784 3776 10848 3780
rect 10864 3836 10928 3840
rect 10864 3780 10868 3836
rect 10868 3780 10924 3836
rect 10924 3780 10928 3836
rect 10864 3776 10928 3780
rect 10944 3836 11008 3840
rect 10944 3780 10948 3836
rect 10948 3780 11004 3836
rect 11004 3780 11008 3836
rect 10944 3776 11008 3780
rect 11024 3836 11088 3840
rect 11024 3780 11028 3836
rect 11028 3780 11084 3836
rect 11084 3780 11088 3836
rect 11024 3776 11088 3780
rect 14717 3836 14781 3840
rect 14717 3780 14721 3836
rect 14721 3780 14777 3836
rect 14777 3780 14781 3836
rect 14717 3776 14781 3780
rect 14797 3836 14861 3840
rect 14797 3780 14801 3836
rect 14801 3780 14857 3836
rect 14857 3780 14861 3836
rect 14797 3776 14861 3780
rect 14877 3836 14941 3840
rect 14877 3780 14881 3836
rect 14881 3780 14937 3836
rect 14937 3780 14941 3836
rect 14877 3776 14941 3780
rect 14957 3836 15021 3840
rect 14957 3780 14961 3836
rect 14961 3780 15017 3836
rect 15017 3780 15021 3836
rect 14957 3776 15021 3780
rect 4884 3292 4948 3296
rect 4884 3236 4888 3292
rect 4888 3236 4944 3292
rect 4944 3236 4948 3292
rect 4884 3232 4948 3236
rect 4964 3292 5028 3296
rect 4964 3236 4968 3292
rect 4968 3236 5024 3292
rect 5024 3236 5028 3292
rect 4964 3232 5028 3236
rect 5044 3292 5108 3296
rect 5044 3236 5048 3292
rect 5048 3236 5104 3292
rect 5104 3236 5108 3292
rect 5044 3232 5108 3236
rect 5124 3292 5188 3296
rect 5124 3236 5128 3292
rect 5128 3236 5184 3292
rect 5184 3236 5188 3292
rect 5124 3232 5188 3236
rect 8817 3292 8881 3296
rect 8817 3236 8821 3292
rect 8821 3236 8877 3292
rect 8877 3236 8881 3292
rect 8817 3232 8881 3236
rect 8897 3292 8961 3296
rect 8897 3236 8901 3292
rect 8901 3236 8957 3292
rect 8957 3236 8961 3292
rect 8897 3232 8961 3236
rect 8977 3292 9041 3296
rect 8977 3236 8981 3292
rect 8981 3236 9037 3292
rect 9037 3236 9041 3292
rect 8977 3232 9041 3236
rect 9057 3292 9121 3296
rect 9057 3236 9061 3292
rect 9061 3236 9117 3292
rect 9117 3236 9121 3292
rect 9057 3232 9121 3236
rect 12750 3292 12814 3296
rect 12750 3236 12754 3292
rect 12754 3236 12810 3292
rect 12810 3236 12814 3292
rect 12750 3232 12814 3236
rect 12830 3292 12894 3296
rect 12830 3236 12834 3292
rect 12834 3236 12890 3292
rect 12890 3236 12894 3292
rect 12830 3232 12894 3236
rect 12910 3292 12974 3296
rect 12910 3236 12914 3292
rect 12914 3236 12970 3292
rect 12970 3236 12974 3292
rect 12910 3232 12974 3236
rect 12990 3292 13054 3296
rect 12990 3236 12994 3292
rect 12994 3236 13050 3292
rect 13050 3236 13054 3292
rect 12990 3232 13054 3236
rect 16683 3292 16747 3296
rect 16683 3236 16687 3292
rect 16687 3236 16743 3292
rect 16743 3236 16747 3292
rect 16683 3232 16747 3236
rect 16763 3292 16827 3296
rect 16763 3236 16767 3292
rect 16767 3236 16823 3292
rect 16823 3236 16827 3292
rect 16763 3232 16827 3236
rect 16843 3292 16907 3296
rect 16843 3236 16847 3292
rect 16847 3236 16903 3292
rect 16903 3236 16907 3292
rect 16843 3232 16907 3236
rect 16923 3292 16987 3296
rect 16923 3236 16927 3292
rect 16927 3236 16983 3292
rect 16983 3236 16987 3292
rect 16923 3232 16987 3236
rect 2918 2748 2982 2752
rect 2918 2692 2922 2748
rect 2922 2692 2978 2748
rect 2978 2692 2982 2748
rect 2918 2688 2982 2692
rect 2998 2748 3062 2752
rect 2998 2692 3002 2748
rect 3002 2692 3058 2748
rect 3058 2692 3062 2748
rect 2998 2688 3062 2692
rect 3078 2748 3142 2752
rect 3078 2692 3082 2748
rect 3082 2692 3138 2748
rect 3138 2692 3142 2748
rect 3078 2688 3142 2692
rect 3158 2748 3222 2752
rect 3158 2692 3162 2748
rect 3162 2692 3218 2748
rect 3218 2692 3222 2748
rect 3158 2688 3222 2692
rect 6851 2748 6915 2752
rect 6851 2692 6855 2748
rect 6855 2692 6911 2748
rect 6911 2692 6915 2748
rect 6851 2688 6915 2692
rect 6931 2748 6995 2752
rect 6931 2692 6935 2748
rect 6935 2692 6991 2748
rect 6991 2692 6995 2748
rect 6931 2688 6995 2692
rect 7011 2748 7075 2752
rect 7011 2692 7015 2748
rect 7015 2692 7071 2748
rect 7071 2692 7075 2748
rect 7011 2688 7075 2692
rect 7091 2748 7155 2752
rect 7091 2692 7095 2748
rect 7095 2692 7151 2748
rect 7151 2692 7155 2748
rect 7091 2688 7155 2692
rect 10784 2748 10848 2752
rect 10784 2692 10788 2748
rect 10788 2692 10844 2748
rect 10844 2692 10848 2748
rect 10784 2688 10848 2692
rect 10864 2748 10928 2752
rect 10864 2692 10868 2748
rect 10868 2692 10924 2748
rect 10924 2692 10928 2748
rect 10864 2688 10928 2692
rect 10944 2748 11008 2752
rect 10944 2692 10948 2748
rect 10948 2692 11004 2748
rect 11004 2692 11008 2748
rect 10944 2688 11008 2692
rect 11024 2748 11088 2752
rect 11024 2692 11028 2748
rect 11028 2692 11084 2748
rect 11084 2692 11088 2748
rect 11024 2688 11088 2692
rect 14717 2748 14781 2752
rect 14717 2692 14721 2748
rect 14721 2692 14777 2748
rect 14777 2692 14781 2748
rect 14717 2688 14781 2692
rect 14797 2748 14861 2752
rect 14797 2692 14801 2748
rect 14801 2692 14857 2748
rect 14857 2692 14861 2748
rect 14797 2688 14861 2692
rect 14877 2748 14941 2752
rect 14877 2692 14881 2748
rect 14881 2692 14937 2748
rect 14937 2692 14941 2748
rect 14877 2688 14941 2692
rect 14957 2748 15021 2752
rect 14957 2692 14961 2748
rect 14961 2692 15017 2748
rect 15017 2692 15021 2748
rect 14957 2688 15021 2692
rect 4884 2204 4948 2208
rect 4884 2148 4888 2204
rect 4888 2148 4944 2204
rect 4944 2148 4948 2204
rect 4884 2144 4948 2148
rect 4964 2204 5028 2208
rect 4964 2148 4968 2204
rect 4968 2148 5024 2204
rect 5024 2148 5028 2204
rect 4964 2144 5028 2148
rect 5044 2204 5108 2208
rect 5044 2148 5048 2204
rect 5048 2148 5104 2204
rect 5104 2148 5108 2204
rect 5044 2144 5108 2148
rect 5124 2204 5188 2208
rect 5124 2148 5128 2204
rect 5128 2148 5184 2204
rect 5184 2148 5188 2204
rect 5124 2144 5188 2148
rect 8817 2204 8881 2208
rect 8817 2148 8821 2204
rect 8821 2148 8877 2204
rect 8877 2148 8881 2204
rect 8817 2144 8881 2148
rect 8897 2204 8961 2208
rect 8897 2148 8901 2204
rect 8901 2148 8957 2204
rect 8957 2148 8961 2204
rect 8897 2144 8961 2148
rect 8977 2204 9041 2208
rect 8977 2148 8981 2204
rect 8981 2148 9037 2204
rect 9037 2148 9041 2204
rect 8977 2144 9041 2148
rect 9057 2204 9121 2208
rect 9057 2148 9061 2204
rect 9061 2148 9117 2204
rect 9117 2148 9121 2204
rect 9057 2144 9121 2148
rect 12750 2204 12814 2208
rect 12750 2148 12754 2204
rect 12754 2148 12810 2204
rect 12810 2148 12814 2204
rect 12750 2144 12814 2148
rect 12830 2204 12894 2208
rect 12830 2148 12834 2204
rect 12834 2148 12890 2204
rect 12890 2148 12894 2204
rect 12830 2144 12894 2148
rect 12910 2204 12974 2208
rect 12910 2148 12914 2204
rect 12914 2148 12970 2204
rect 12970 2148 12974 2204
rect 12910 2144 12974 2148
rect 12990 2204 13054 2208
rect 12990 2148 12994 2204
rect 12994 2148 13050 2204
rect 13050 2148 13054 2204
rect 12990 2144 13054 2148
rect 16683 2204 16747 2208
rect 16683 2148 16687 2204
rect 16687 2148 16743 2204
rect 16743 2148 16747 2204
rect 16683 2144 16747 2148
rect 16763 2204 16827 2208
rect 16763 2148 16767 2204
rect 16767 2148 16823 2204
rect 16823 2148 16827 2204
rect 16763 2144 16827 2148
rect 16843 2204 16907 2208
rect 16843 2148 16847 2204
rect 16847 2148 16903 2204
rect 16903 2148 16907 2204
rect 16843 2144 16907 2148
rect 16923 2204 16987 2208
rect 16923 2148 16927 2204
rect 16927 2148 16983 2204
rect 16983 2148 16987 2204
rect 16923 2144 16987 2148
<< metal4 >>
rect 2910 15808 3230 15824
rect 2910 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3230 15808
rect 2910 14720 3230 15744
rect 2910 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3230 14720
rect 2910 13632 3230 14656
rect 2910 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3230 13632
rect 2910 12544 3230 13568
rect 2910 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3230 12544
rect 2910 11456 3230 12480
rect 2910 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3230 11456
rect 2910 10368 3230 11392
rect 2910 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3230 10368
rect 2910 9280 3230 10304
rect 2910 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3230 9280
rect 2910 8192 3230 9216
rect 2910 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3230 8192
rect 2910 7104 3230 8128
rect 2910 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3230 7104
rect 2910 6016 3230 7040
rect 2910 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3230 6016
rect 2910 4928 3230 5952
rect 2910 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3230 4928
rect 2910 3840 3230 4864
rect 2910 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3230 3840
rect 2910 2752 3230 3776
rect 2910 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3230 2752
rect 2910 2128 3230 2688
rect 4876 15264 5196 15824
rect 4876 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5196 15264
rect 4876 14176 5196 15200
rect 4876 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5196 14176
rect 4876 13088 5196 14112
rect 4876 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5196 13088
rect 4876 12000 5196 13024
rect 4876 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5196 12000
rect 4876 10912 5196 11936
rect 4876 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5196 10912
rect 4876 9824 5196 10848
rect 4876 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5196 9824
rect 4876 8736 5196 9760
rect 4876 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5196 8736
rect 4876 7648 5196 8672
rect 4876 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5196 7648
rect 4876 6560 5196 7584
rect 4876 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5196 6560
rect 4876 5472 5196 6496
rect 4876 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5196 5472
rect 4876 4384 5196 5408
rect 4876 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5196 4384
rect 4876 3296 5196 4320
rect 4876 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5196 3296
rect 4876 2208 5196 3232
rect 4876 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5196 2208
rect 4876 2128 5196 2144
rect 6843 15808 7163 15824
rect 6843 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7163 15808
rect 6843 14720 7163 15744
rect 6843 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7163 14720
rect 6843 13632 7163 14656
rect 6843 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7163 13632
rect 6843 12544 7163 13568
rect 6843 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7163 12544
rect 6843 11456 7163 12480
rect 6843 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7163 11456
rect 6843 10368 7163 11392
rect 6843 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7163 10368
rect 6843 9280 7163 10304
rect 6843 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7163 9280
rect 6843 8192 7163 9216
rect 6843 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7163 8192
rect 6843 7104 7163 8128
rect 6843 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7163 7104
rect 6843 6016 7163 7040
rect 6843 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7163 6016
rect 6843 4928 7163 5952
rect 6843 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7163 4928
rect 6843 3840 7163 4864
rect 6843 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7163 3840
rect 6843 2752 7163 3776
rect 6843 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7163 2752
rect 6843 2128 7163 2688
rect 8809 15264 9129 15824
rect 8809 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9129 15264
rect 8809 14176 9129 15200
rect 8809 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9129 14176
rect 8809 13088 9129 14112
rect 8809 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9129 13088
rect 8809 12000 9129 13024
rect 8809 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9129 12000
rect 8809 10912 9129 11936
rect 8809 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9129 10912
rect 8809 9824 9129 10848
rect 8809 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9129 9824
rect 8809 8736 9129 9760
rect 8809 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9129 8736
rect 8809 7648 9129 8672
rect 8809 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9129 7648
rect 8809 6560 9129 7584
rect 8809 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9129 6560
rect 8809 5472 9129 6496
rect 8809 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9129 5472
rect 8809 4384 9129 5408
rect 8809 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9129 4384
rect 8809 3296 9129 4320
rect 8809 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9129 3296
rect 8809 2208 9129 3232
rect 8809 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9129 2208
rect 8809 2128 9129 2144
rect 10776 15808 11096 15824
rect 10776 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11096 15808
rect 10776 14720 11096 15744
rect 10776 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11096 14720
rect 10776 13632 11096 14656
rect 10776 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11096 13632
rect 10776 12544 11096 13568
rect 10776 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11096 12544
rect 10776 11456 11096 12480
rect 10776 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11096 11456
rect 10776 10368 11096 11392
rect 10776 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11096 10368
rect 10776 9280 11096 10304
rect 10776 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11096 9280
rect 10776 8192 11096 9216
rect 10776 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11096 8192
rect 10776 7104 11096 8128
rect 10776 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11096 7104
rect 10776 6016 11096 7040
rect 10776 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11096 6016
rect 10776 4928 11096 5952
rect 10776 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11096 4928
rect 10776 3840 11096 4864
rect 10776 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11096 3840
rect 10776 2752 11096 3776
rect 10776 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11096 2752
rect 10776 2128 11096 2688
rect 12742 15264 13062 15824
rect 12742 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13062 15264
rect 12742 14176 13062 15200
rect 12742 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13062 14176
rect 12742 13088 13062 14112
rect 12742 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13062 13088
rect 12742 12000 13062 13024
rect 12742 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13062 12000
rect 12742 10912 13062 11936
rect 12742 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13062 10912
rect 12742 9824 13062 10848
rect 12742 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13062 9824
rect 12742 8736 13062 9760
rect 12742 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13062 8736
rect 12742 7648 13062 8672
rect 12742 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13062 7648
rect 12742 6560 13062 7584
rect 12742 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13062 6560
rect 12742 5472 13062 6496
rect 12742 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13062 5472
rect 12742 4384 13062 5408
rect 12742 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13062 4384
rect 12742 3296 13062 4320
rect 12742 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13062 3296
rect 12742 2208 13062 3232
rect 12742 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13062 2208
rect 12742 2128 13062 2144
rect 14709 15808 15029 15824
rect 14709 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15029 15808
rect 14709 14720 15029 15744
rect 14709 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15029 14720
rect 14709 13632 15029 14656
rect 14709 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15029 13632
rect 14709 12544 15029 13568
rect 14709 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15029 12544
rect 14709 11456 15029 12480
rect 14709 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15029 11456
rect 14709 10368 15029 11392
rect 14709 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15029 10368
rect 14709 9280 15029 10304
rect 14709 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15029 9280
rect 14709 8192 15029 9216
rect 14709 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15029 8192
rect 14709 7104 15029 8128
rect 14709 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15029 7104
rect 14709 6016 15029 7040
rect 14709 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15029 6016
rect 14709 4928 15029 5952
rect 14709 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15029 4928
rect 14709 3840 15029 4864
rect 14709 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15029 3840
rect 14709 2752 15029 3776
rect 14709 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15029 2752
rect 14709 2128 15029 2688
rect 16675 15264 16995 15824
rect 16675 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16995 15264
rect 16675 14176 16995 15200
rect 16675 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16995 14176
rect 16675 13088 16995 14112
rect 16675 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16995 13088
rect 16675 12000 16995 13024
rect 16675 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16995 12000
rect 16675 10912 16995 11936
rect 16675 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16995 10912
rect 16675 9824 16995 10848
rect 16675 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16995 9824
rect 16675 8736 16995 9760
rect 16675 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16995 8736
rect 16675 7648 16995 8672
rect 16675 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16995 7648
rect 16675 6560 16995 7584
rect 16675 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16995 6560
rect 16675 5472 16995 6496
rect 16675 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16995 5472
rect 16675 4384 16995 5408
rect 16675 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16995 4384
rect 16675 3296 16995 4320
rect 16675 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16995 3296
rect 16675 2208 16995 3232
rect 16675 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16995 2208
rect 16675 2128 16995 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_spi_clk_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1673029049
transform -1 0 2392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1673029049
transform -1 0 2944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1673029049
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1673029049
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1673029049
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1673029049
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1673029049
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1673029049
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1673029049
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1673029049
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1673029049
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1673029049
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1673029049
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1673029049
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1673029049
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1673029049
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1673029049
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1673029049
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1673029049
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1673029049
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1673029049
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1673029049
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1673029049
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1673029049
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1673029049
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1673029049
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1673029049
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1673029049
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1673029049
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1673029049
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1673029049
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1673029049
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1673029049
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1673029049
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1673029049
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1673029049
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1673029049
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1673029049
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1673029049
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1673029049
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1673029049
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1673029049
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1673029049
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1673029049
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1673029049
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1673029049
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1673029049
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1673029049
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1673029049
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1673029049
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_165
timestamp 1673029049
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1673029049
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1673029049
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1673029049
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1673029049
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1673029049
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1673029049
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1673029049
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1673029049
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1673029049
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1673029049
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1673029049
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1673029049
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1673029049
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1673029049
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1673029049
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1673029049
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1673029049
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1673029049
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1673029049
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1673029049
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1673029049
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1673029049
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1673029049
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1673029049
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1673029049
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1673029049
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1673029049
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1673029049
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1673029049
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1673029049
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1673029049
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1673029049
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1673029049
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1673029049
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1673029049
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 1673029049
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1673029049
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1673029049
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1673029049
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1673029049
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1673029049
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1673029049
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1673029049
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1673029049
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1673029049
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1673029049
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1673029049
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1673029049
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1673029049
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1673029049
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1673029049
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1673029049
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1673029049
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1673029049
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1673029049
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1673029049
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1673029049
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1673029049
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1673029049
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1673029049
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1673029049
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1673029049
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1673029049
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1673029049
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1673029049
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1673029049
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1673029049
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1673029049
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1673029049
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1673029049
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1673029049
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 1673029049
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1673029049
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1673029049
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1673029049
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1673029049
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1673029049
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1673029049
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1673029049
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1673029049
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1673029049
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1673029049
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1673029049
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1673029049
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1673029049
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1673029049
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1673029049
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1673029049
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1673029049
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1673029049
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1673029049
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1673029049
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_14
timestamp 1673029049
transform 1 0 2392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1673029049
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1673029049
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1673029049
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1673029049
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1673029049
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1673029049
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1673029049
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1673029049
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1673029049
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1673029049
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1673029049
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1673029049
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1673029049
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1673029049
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1673029049
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp 1673029049
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1673029049
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1673029049
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1673029049
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1673029049
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1673029049
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1673029049
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1673029049
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1673029049
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1673029049
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1673029049
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1673029049
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1673029049
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1673029049
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1673029049
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1673029049
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1673029049
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1673029049
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1673029049
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1673029049
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1673029049
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1673029049
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1673029049
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1673029049
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1673029049
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1673029049
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1673029049
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1673029049
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1673029049
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1673029049
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1673029049
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1673029049
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1673029049
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1673029049
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1673029049
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1673029049
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp 1673029049
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1673029049
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1673029049
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1673029049
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1673029049
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1673029049
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1673029049
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1673029049
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1673029049
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1673029049
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1673029049
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1673029049
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1673029049
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1673029049
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1673029049
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1673029049
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1673029049
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1673029049
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1673029049
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1673029049
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1673029049
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1673029049
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1673029049
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1673029049
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1673029049
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1673029049
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1673029049
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1673029049
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1673029049
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1673029049
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1673029049
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1673029049
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1673029049
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1673029049
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1673029049
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1673029049
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1673029049
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1673029049
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_165
timestamp 1673029049
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_11
timestamp 1673029049
transform 1 0 2116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1673029049
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_23
timestamp 1673029049
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_33
timestamp 1673029049
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1673029049
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1673029049
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1673029049
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1673029049
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1673029049
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1673029049
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1673029049
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1673029049
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1673029049
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1673029049
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1673029049
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1673029049
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1673029049
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1673029049
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1673029049
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_9
timestamp 1673029049
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1673029049
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1673029049
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1673029049
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_38
timestamp 1673029049
transform 1 0 4600 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_50
timestamp 1673029049
transform 1 0 5704 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_62
timestamp 1673029049
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_72
timestamp 1673029049
transform 1 0 7728 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1673029049
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1673029049
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1673029049
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1673029049
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1673029049
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1673029049
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1673029049
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1673029049
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_165
timestamp 1673029049
transform 1 0 16284 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1673029049
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_14
timestamp 1673029049
transform 1 0 2392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_20
timestamp 1673029049
transform 1 0 2944 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_34
timestamp 1673029049
transform 1 0 4232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1673029049
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1673029049
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1673029049
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_65
timestamp 1673029049
transform 1 0 7084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_77
timestamp 1673029049
transform 1 0 8188 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_89
timestamp 1673029049
transform 1 0 9292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp 1673029049
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1673029049
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1673029049
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1673029049
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1673029049
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1673029049
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1673029049
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1673029049
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1673029049
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_9
timestamp 1673029049
transform 1 0 1932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_15
timestamp 1673029049
transform 1 0 2484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_19
timestamp 1673029049
transform 1 0 2852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1673029049
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1673029049
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_44
timestamp 1673029049
transform 1 0 5152 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_54
timestamp 1673029049
transform 1 0 6072 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_66
timestamp 1673029049
transform 1 0 7176 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 1673029049
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1673029049
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1673029049
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1673029049
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1673029049
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1673029049
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1673029049
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1673029049
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1673029049
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_165
timestamp 1673029049
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1673029049
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_17
timestamp 1673029049
transform 1 0 2668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_33
timestamp 1673029049
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_41
timestamp 1673029049
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1673029049
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1673029049
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1673029049
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_63
timestamp 1673029049
transform 1 0 6900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_75
timestamp 1673029049
transform 1 0 8004 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1673029049
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1673029049
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1673029049
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1673029049
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1673029049
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1673029049
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1673029049
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1673029049
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1673029049
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1673029049
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1673029049
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1673029049
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1673029049
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1673029049
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1673029049
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_62
timestamp 1673029049
transform 1 0 6808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1673029049
transform 1 0 7912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1673029049
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1673029049
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1673029049
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1673029049
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1673029049
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1673029049
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1673029049
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1673029049
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1673029049
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_165
timestamp 1673029049
transform 1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1673029049
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1673029049
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_36
timestamp 1673029049
transform 1 0 4416 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1673029049
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1673029049
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1673029049
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_66
timestamp 1673029049
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_78
timestamp 1673029049
transform 1 0 8280 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_90
timestamp 1673029049
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1673029049
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1673029049
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1673029049
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1673029049
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1673029049
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1673029049
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1673029049
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1673029049
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1673029049
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1673029049
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1673029049
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_51
timestamp 1673029049
transform 1 0 5796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1673029049
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_62
timestamp 1673029049
transform 1 0 6808 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_70
timestamp 1673029049
transform 1 0 7544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1673029049
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1673029049
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1673029049
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1673029049
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1673029049
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1673029049
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1673029049
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1673029049
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1673029049
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1673029049
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1673029049
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_13
timestamp 1673029049
transform 1 0 2300 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_21
timestamp 1673029049
transform 1 0 3036 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_43
timestamp 1673029049
transform 1 0 5060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_47
timestamp 1673029049
transform 1 0 5428 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1673029049
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1673029049
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1673029049
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_68
timestamp 1673029049
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_80
timestamp 1673029049
transform 1 0 8464 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_92
timestamp 1673029049
transform 1 0 9568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1673029049
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1673029049
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1673029049
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1673029049
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1673029049
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1673029049
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1673029049
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1673029049
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1673029049
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1673029049
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1673029049
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1673029049
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1673029049
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1673029049
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1673029049
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1673029049
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1673029049
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1673029049
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1673029049
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1673029049
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1673029049
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1673029049
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1673029049
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_17
timestamp 1673029049
transform 1 0 2668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1673029049
transform 1 0 5152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1673029049
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1673029049
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_61
timestamp 1673029049
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_65
timestamp 1673029049
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_78
timestamp 1673029049
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_90
timestamp 1673029049
transform 1 0 9384 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1673029049
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1673029049
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1673029049
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1673029049
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1673029049
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1673029049
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1673029049
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1673029049
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1673029049
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_10
timestamp 1673029049
transform 1 0 2024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_17
timestamp 1673029049
transform 1 0 2668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1673029049
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1673029049
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1673029049
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1673029049
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_54
timestamp 1673029049
transform 1 0 6072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_57
timestamp 1673029049
transform 1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_62
timestamp 1673029049
transform 1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1673029049
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1673029049
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1673029049
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1673029049
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1673029049
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_106
timestamp 1673029049
transform 1 0 10856 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_113
timestamp 1673029049
transform 1 0 11500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_125
timestamp 1673029049
transform 1 0 12604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1673029049
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1673029049
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_153
timestamp 1673029049
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_161
timestamp 1673029049
transform 1 0 15916 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_166
timestamp 1673029049
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1673029049
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1673029049
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1673029049
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1673029049
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1673029049
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1673029049
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1673029049
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1673029049
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1673029049
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1673029049
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1673029049
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1673029049
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1673029049
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1673029049
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1673029049
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1673029049
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1673029049
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1673029049
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1673029049
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1673029049
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1673029049
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1673029049
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1673029049
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1673029049
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1673029049
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1673029049
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1673029049
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1673029049
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1673029049
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1673029049
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1673029049
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1673029049
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1673029049
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1673029049
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1673029049
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1673029049
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1673029049
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1673029049
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1673029049
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1673029049
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1673029049
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1673029049
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1673029049
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1673029049
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1673029049
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1673029049
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1673029049
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1673029049
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1673029049
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1673029049
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1673029049
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1673029049
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1673029049
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1673029049
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1673029049
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1673029049
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1673029049
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1673029049
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1673029049
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1673029049
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1673029049
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1673029049
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1673029049
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1673029049
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1673029049
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1673029049
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1673029049
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1673029049
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1673029049
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1673029049
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1673029049
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1673029049
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1673029049
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1673029049
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1673029049
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1673029049
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1673029049
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1673029049
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1673029049
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1673029049
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1673029049
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1673029049
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1673029049
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1673029049
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1673029049
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1673029049
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1673029049
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1673029049
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1673029049
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1673029049
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1673029049
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1673029049
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _32_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _33_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6900 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _34_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _35_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 7360 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _36_
timestamp 1673029049
transform -1 0 6072 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _37_
timestamp 1673029049
transform -1 0 4140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _38_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _39_
timestamp 1673029049
transform -1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _40_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _41_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6348 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1673029049
transform -1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _43_
timestamp 1673029049
transform -1 0 7176 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _44_
timestamp 1673029049
transform -1 0 6072 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _45_
timestamp 1673029049
transform 1 0 1932 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _46_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3680 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1673029049
transform 1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1673029049
transform -1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1673029049
transform -1 0 2852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _50_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3404 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _51_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 7728 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _52_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5520 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _53_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _54_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _55_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 2300 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _56_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _57_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3956 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1673029049
transform -1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1673029049
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1673029049
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _61_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _62_
timestamp 1673029049
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _63_
timestamp 1673029049
transform 1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _64_
timestamp 1673029049
transform -1 0 3312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _65_
timestamp 1673029049
transform 1 0 6164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _66_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _67_
timestamp 1673029049
transform 1 0 7176 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _68_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3128 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _69_
timestamp 1673029049
transform 1 0 3956 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _70_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3956 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _71_
timestamp 1673029049
transform 1 0 1564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _72_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3036 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dlxtn_1  _73_
timestamp 1673029049
transform -1 0 2668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _74_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 5152 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _75_
timestamp 1673029049
transform -1 0 2668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _76_
timestamp 1673029049
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _77_
timestamp 1673029049
transform -1 0 6072 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_spi_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 3496 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_spi_clk
timestamp 1673029049
transform -1 0 3404 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_spi_clk
timestamp 1673029049
transform 1 0 2576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1673029049
transform -1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1673029049
transform -1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1673029049
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1673029049
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1673029049
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1673029049
transform -1 0 2024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1673029049
transform 1 0 1564 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 4526 17200 4582 18000 0 FreeSans 224 90 0 0 reg_addr[0]
port 0 nsew signal tristate
flabel metal2 s 7470 17200 7526 18000 0 FreeSans 224 90 0 0 reg_addr[1]
port 1 nsew signal tristate
flabel metal2 s 10414 17200 10470 18000 0 FreeSans 224 90 0 0 reg_addr[2]
port 2 nsew signal tristate
flabel metal2 s 13358 17200 13414 18000 0 FreeSans 224 90 0 0 reg_bus
port 3 nsew signal bidirectional
flabel metal2 s 16302 17200 16358 18000 0 FreeSans 224 90 0 0 reg_clk
port 4 nsew signal tristate
flabel metal2 s 1582 17200 1638 18000 0 FreeSans 224 90 0 0 reg_dir
port 5 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 spi_clk
port 6 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 spi_miso
port 7 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 spi_mosi
port 8 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 spi_sel
port 9 nsew signal input
flabel metal4 s 2910 2128 3230 15824 0 FreeSans 1920 90 0 0 vcc
port 10 nsew power bidirectional
flabel metal4 s 6843 2128 7163 15824 0 FreeSans 1920 90 0 0 vcc
port 10 nsew power bidirectional
flabel metal4 s 10776 2128 11096 15824 0 FreeSans 1920 90 0 0 vcc
port 10 nsew power bidirectional
flabel metal4 s 14709 2128 15029 15824 0 FreeSans 1920 90 0 0 vcc
port 10 nsew power bidirectional
flabel metal4 s 4876 2128 5196 15824 0 FreeSans 1920 90 0 0 vss
port 11 nsew ground bidirectional
flabel metal4 s 8809 2128 9129 15824 0 FreeSans 1920 90 0 0 vss
port 11 nsew ground bidirectional
flabel metal4 s 12742 2128 13062 15824 0 FreeSans 1920 90 0 0 vss
port 11 nsew ground bidirectional
flabel metal4 s 16675 2128 16995 15824 0 FreeSans 1920 90 0 0 vss
port 11 nsew ground bidirectional
rlabel metal1 8970 15776 8970 15776 0 vcc
rlabel via1 9049 15232 9049 15232 0 vss
rlabel metal1 2346 15062 2346 15062 0 _00_
rlabel metal1 8878 11764 8878 11764 0 _01_
rlabel metal2 3450 12852 3450 12852 0 _02_
rlabel metal1 5704 11254 5704 11254 0 _03_
rlabel metal1 4692 11866 4692 11866 0 _04_
rlabel metal1 2346 9146 2346 9146 0 _05_
rlabel metal1 6118 10778 6118 10778 0 _06_
rlabel metal1 3450 11254 3450 11254 0 _07_
rlabel metal2 8602 11900 8602 11900 0 _08_
rlabel metal2 6026 14722 6026 14722 0 _09_
rlabel metal1 6302 14348 6302 14348 0 _10_
rlabel metal1 6624 14926 6624 14926 0 _11_
rlabel metal1 2990 10234 2990 10234 0 _12_
rlabel metal2 3726 14824 3726 14824 0 _13_
rlabel metal2 3726 13056 3726 13056 0 _14_
rlabel metal1 3181 13226 3181 13226 0 _15_
rlabel metal2 6302 14280 6302 14280 0 _16_
rlabel via2 5658 13923 5658 13923 0 _17_
rlabel metal1 7636 13498 7636 13498 0 _18_
rlabel metal1 5380 11730 5380 11730 0 _19_
rlabel metal2 1886 9146 1886 9146 0 _20_
rlabel metal1 5980 12614 5980 12614 0 _21_
rlabel metal1 7544 12206 7544 12206 0 _22_
rlabel metal1 6072 12954 6072 12954 0 _23_
rlabel metal1 3036 10642 3036 10642 0 _24_
rlabel metal1 4508 10778 4508 10778 0 _25_
rlabel metal2 2438 10268 2438 10268 0 _26_
rlabel metal1 5750 11084 5750 11084 0 _27_
rlabel metal2 5290 11968 5290 11968 0 _28_
rlabel metal1 1610 13940 1610 13940 0 _29_
rlabel metal2 4554 10438 4554 10438 0 _30_
rlabel metal1 3496 11118 3496 11118 0 _31_
rlabel metal1 2392 12886 2392 12886 0 clknet_0_spi_clk
rlabel metal1 2295 14042 2295 14042 0 clknet_1_0__leaf_spi_clk
rlabel metal1 3956 13294 3956 13294 0 clknet_1_1__leaf_spi_clk
rlabel metal1 1794 6664 1794 6664 0 net1
rlabel metal2 1886 12036 1886 12036 0 net2
rlabel metal1 4784 15470 4784 15470 0 net3
rlabel metal1 7452 14586 7452 14586 0 net4
rlabel metal1 8280 15130 8280 15130 0 net5
rlabel metal1 1840 15130 1840 15130 0 net6
rlabel metal1 1978 15538 1978 15538 0 net7
rlabel metal2 1610 6970 1610 6970 0 net8
rlabel via1 4646 12415 4646 12415 0 next_state\[0\]
rlabel metal1 3082 11322 3082 11322 0 next_state\[1\]
rlabel metal1 6578 11662 6578 11662 0 pres_state\[0\]
rlabel metal1 2208 10642 2208 10642 0 pres_state\[1\]
rlabel metal1 4462 15674 4462 15674 0 reg_addr[0]
rlabel metal1 7636 15674 7636 15674 0 reg_addr[1]
rlabel metal2 10718 16507 10718 16507 0 reg_addr[2]
rlabel metal1 2898 11730 2898 11730 0 reg_bus
rlabel metal2 16277 17340 16277 17340 0 reg_clk
rlabel metal1 1702 15674 1702 15674 0 reg_dir
rlabel metal1 3128 14382 3128 14382 0 spi_clk
rlabel metal3 1234 2244 1234 2244 0 spi_miso
rlabel metal1 1564 6766 1564 6766 0 spi_mosi
rlabel metal2 1702 11169 1702 11169 0 spi_sel
rlabel metal1 5428 12206 5428 12206 0 t\[0\]
rlabel metal1 5612 12274 5612 12274 0 t\[1\]
rlabel metal1 5842 12274 5842 12274 0 t\[2\]
<< properties >>
string FIXED_BBOX 0 0 18000 18000
<< end >>
