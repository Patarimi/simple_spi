VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spi_register
  CLASS BLOCK ;
  FOREIGN spi_register ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END reg_addr[2]
  PIN reg_bus
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END reg_bus
  PIN reg_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END reg_clk
  PIN reg_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 116.000 8.650 120.000 ;
    END
  END reg_data[0]
  PIN reg_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 116.000 23.370 120.000 ;
    END
  END reg_data[1]
  PIN reg_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 116.000 38.090 120.000 ;
    END
  END reg_data[2]
  PIN reg_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 116.000 52.810 120.000 ;
    END
  END reg_data[3]
  PIN reg_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 116.000 67.530 120.000 ;
    END
  END reg_data[4]
  PIN reg_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 116.000 82.250 120.000 ;
    END
  END reg_data[5]
  PIN reg_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 116.000 96.970 120.000 ;
    END
  END reg_data[6]
  PIN reg_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 116.000 111.690 120.000 ;
    END
  END reg_data[7]
  PIN reg_dir
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END reg_dir
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.290 10.640 19.890 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.430 10.640 47.030 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.570 10.640 74.170 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.710 10.640 101.310 109.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 31.860 10.640 33.460 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.000 10.640 60.600 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.140 10.640 87.740 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.280 10.640 114.880 109.040 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 104.665 114.270 107.495 ;
        RECT 5.330 99.225 114.270 102.055 ;
        RECT 5.330 93.785 114.270 96.615 ;
        RECT 5.330 88.345 114.270 91.175 ;
        RECT 5.330 82.905 114.270 85.735 ;
        RECT 5.330 77.465 114.270 80.295 ;
        RECT 5.330 72.025 114.270 74.855 ;
        RECT 5.330 66.585 114.270 69.415 ;
        RECT 5.330 61.145 114.270 63.975 ;
        RECT 5.330 55.705 114.270 58.535 ;
        RECT 5.330 50.265 114.270 53.095 ;
        RECT 5.330 44.825 114.270 47.655 ;
        RECT 5.330 39.385 114.270 42.215 ;
        RECT 5.330 33.945 114.270 36.775 ;
        RECT 5.330 28.505 114.270 31.335 ;
        RECT 5.330 23.065 114.270 25.895 ;
        RECT 5.330 17.625 114.270 20.455 ;
        RECT 5.330 12.185 114.270 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 5.520 10.640 114.880 109.040 ;
      LAYER met2 ;
        RECT 8.930 115.720 22.810 116.690 ;
        RECT 23.650 115.720 37.530 116.690 ;
        RECT 38.370 115.720 52.250 116.690 ;
        RECT 53.090 115.720 66.970 116.690 ;
        RECT 67.810 115.720 81.690 116.690 ;
        RECT 82.530 115.720 96.410 116.690 ;
        RECT 97.250 115.720 111.130 116.690 ;
        RECT 111.970 115.720 114.850 116.690 ;
        RECT 8.650 4.280 114.850 115.720 ;
        RECT 8.650 4.000 9.930 4.280 ;
        RECT 10.770 4.000 29.710 4.280 ;
        RECT 30.550 4.000 49.490 4.280 ;
        RECT 50.330 4.000 69.270 4.280 ;
        RECT 70.110 4.000 89.050 4.280 ;
        RECT 89.890 4.000 108.830 4.280 ;
        RECT 109.670 4.000 114.850 4.280 ;
      LAYER met3 ;
        RECT 18.300 10.715 114.870 108.965 ;
  END
END spi_register
END LIBRARY

