magic
tech sky130A
magscale 1 2
timestamp 1672930028
<< viali >>
rect 7389 7497 7423 7531
rect 8401 7497 8435 7531
rect 3433 7361 3467 7395
rect 4629 7361 4663 7395
rect 5273 7361 5307 7395
rect 6009 7361 6043 7395
rect 7205 7361 7239 7395
rect 8585 7361 8619 7395
rect 9229 7361 9263 7395
rect 10517 7361 10551 7395
rect 10977 7361 11011 7395
rect 11713 7361 11747 7395
rect 14933 7361 14967 7395
rect 2145 7293 2179 7327
rect 6745 7293 6779 7327
rect 12357 7293 12391 7327
rect 13001 7293 13035 7327
rect 17509 7293 17543 7327
rect 2789 7225 2823 7259
rect 14289 7225 14323 7259
rect 15577 7225 15611 7259
rect 5825 7157 5859 7191
rect 9321 7157 9355 7191
rect 16865 7157 16899 7191
rect 18153 7157 18187 7191
rect 5181 6953 5215 6987
rect 9229 6953 9263 6987
rect 15577 6953 15611 6987
rect 16221 6885 16255 6919
rect 16865 6885 16899 6919
rect 2145 6817 2179 6851
rect 6469 6817 6503 6851
rect 7849 6817 7883 6851
rect 9873 6817 9907 6851
rect 10517 6817 10551 6851
rect 10977 6817 11011 6851
rect 11621 6817 11655 6851
rect 12909 6817 12943 6851
rect 2789 6749 2823 6783
rect 3433 6749 3467 6783
rect 4537 6749 4571 6783
rect 5825 6749 5859 6783
rect 6929 6749 6963 6783
rect 8585 6749 8619 6783
rect 12265 6749 12299 6783
rect 13553 6749 13587 6783
rect 14289 6749 14323 6783
rect 14933 6749 14967 6783
rect 17509 6749 17543 6783
rect 7113 6613 7147 6647
rect 8401 6613 8435 6647
rect 12725 6409 12759 6443
rect 2605 6273 2639 6307
rect 5273 6273 5307 6307
rect 7021 6273 7055 6307
rect 7481 6273 7515 6307
rect 7665 6273 7699 6307
rect 8769 6273 8803 6307
rect 10057 6273 10091 6307
rect 10517 6273 10551 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 13461 6273 13495 6307
rect 14197 6273 14231 6307
rect 14841 6273 14875 6307
rect 16865 6273 16899 6307
rect 3893 6205 3927 6239
rect 4997 6205 5031 6239
rect 13737 6205 13771 6239
rect 16129 6205 16163 6239
rect 1961 6137 1995 6171
rect 6009 6137 6043 6171
rect 7849 6137 7883 6171
rect 9413 6137 9447 6171
rect 15485 6137 15519 6171
rect 3249 6069 3283 6103
rect 4537 6069 4571 6103
rect 11897 6069 11931 6103
rect 12173 6069 12207 6103
rect 4813 5865 4847 5899
rect 6653 5865 6687 5899
rect 7757 5865 7791 5899
rect 8585 5865 8619 5899
rect 10609 5865 10643 5899
rect 13553 5865 13587 5899
rect 15577 5865 15611 5899
rect 7389 5797 7423 5831
rect 10149 5797 10183 5831
rect 14933 5797 14967 5831
rect 3341 5729 3375 5763
rect 11529 5729 11563 5763
rect 14289 5729 14323 5763
rect 1593 5661 1627 5695
rect 3985 5661 4019 5695
rect 4905 5661 4939 5695
rect 5181 5661 5215 5695
rect 5641 5661 5675 5695
rect 5917 5661 5951 5695
rect 9137 5661 9171 5695
rect 9413 5661 9447 5695
rect 11253 5661 11287 5695
rect 1869 5593 1903 5627
rect 4169 5525 4203 5559
rect 4629 5525 4663 5559
rect 7757 5525 7791 5559
rect 7941 5525 7975 5559
rect 13001 5525 13035 5559
rect 5549 5321 5583 5355
rect 7757 5321 7791 5355
rect 12081 5321 12115 5355
rect 12265 5321 12299 5355
rect 12909 5321 12943 5355
rect 1593 5185 1627 5219
rect 3709 5185 3743 5219
rect 4169 5191 4203 5225
rect 4353 5185 4387 5219
rect 5163 5185 5197 5219
rect 5273 5207 5307 5241
rect 5365 5207 5399 5241
rect 6745 5185 6779 5219
rect 7297 5185 7331 5219
rect 7573 5185 7607 5219
rect 8677 5185 8711 5219
rect 9137 5185 9171 5219
rect 9873 5185 9907 5219
rect 11713 5185 11747 5219
rect 12725 5185 12759 5219
rect 13369 5185 13403 5219
rect 14657 5185 14691 5219
rect 15301 5185 15335 5219
rect 2421 5117 2455 5151
rect 3065 5049 3099 5083
rect 7389 5049 7423 5083
rect 7481 5049 7515 5083
rect 1777 4981 1811 5015
rect 4353 4981 4387 5015
rect 4537 4981 4571 5015
rect 12081 4981 12115 5015
rect 13553 4981 13587 5015
rect 5641 4777 5675 4811
rect 6377 4777 6411 4811
rect 9321 4777 9355 4811
rect 12817 4777 12851 4811
rect 13553 4777 13587 4811
rect 4169 4709 4203 4743
rect 4997 4709 5031 4743
rect 1685 4641 1719 4675
rect 10517 4641 10551 4675
rect 6837 4573 6871 4607
rect 9137 4573 9171 4607
rect 9873 4573 9907 4607
rect 12725 4573 12759 4607
rect 13369 4573 13403 4607
rect 1961 4505 1995 4539
rect 4445 4505 4479 4539
rect 5457 4505 5491 4539
rect 7113 4505 7147 4539
rect 10793 4505 10827 4539
rect 3433 4437 3467 4471
rect 3985 4437 4019 4471
rect 5657 4437 5691 4471
rect 5825 4437 5859 4471
rect 8585 4437 8619 4471
rect 10057 4437 10091 4471
rect 12265 4437 12299 4471
rect 7573 4233 7607 4267
rect 8401 4165 8435 4199
rect 2513 4097 2547 4131
rect 3065 4097 3099 4131
rect 3157 4097 3191 4131
rect 3893 4097 3927 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 5549 4097 5583 4131
rect 6561 4097 6595 4131
rect 7389 4097 7423 4131
rect 7665 4097 7699 4131
rect 8125 4097 8159 4131
rect 8217 4097 8251 4131
rect 8861 4097 8895 4131
rect 11805 4097 11839 4131
rect 11897 4097 11931 4131
rect 2329 3961 2363 3995
rect 4077 3961 4111 3995
rect 4721 3961 4755 3995
rect 9045 3961 9079 3995
rect 7205 3893 7239 3927
rect 8125 3893 8159 3927
rect 2329 3689 2363 3723
rect 3065 3689 3099 3723
rect 4997 3689 5031 3723
rect 5733 3689 5767 3723
rect 6653 3689 6687 3723
rect 7297 3689 7331 3723
rect 8493 3689 8527 3723
rect 7481 3621 7515 3655
rect 2513 3485 2547 3519
rect 3157 3485 3191 3519
rect 6469 3485 6503 3519
rect 8585 3485 8619 3519
rect 7113 3417 7147 3451
rect 7329 3417 7363 3451
rect 5457 3145 5491 3179
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
<< metal1 >>
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 14918 8276 14924 8288
rect 12860 8248 14924 8276
rect 12860 8236 12866 8248
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 8662 8004 8668 8016
rect 5316 7976 8668 8004
rect 5316 7964 5322 7976
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 9214 7936 9220 7948
rect 8628 7908 9220 7936
rect 8628 7896 8634 7908
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 7650 7800 7656 7812
rect 7340 7772 7656 7800
rect 7340 7760 7346 7772
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 7926 7732 7932 7744
rect 4672 7704 7932 7732
rect 4672 7692 4678 7704
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 8846 7732 8852 7744
rect 8444 7704 8852 7732
rect 8444 7692 8450 7704
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 14642 7732 14648 7744
rect 12952 7704 14648 7732
rect 12952 7692 12958 7704
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 1104 7642 18860 7664
rect 1104 7590 3829 7642
rect 3881 7590 3893 7642
rect 3945 7590 3957 7642
rect 4009 7590 4021 7642
rect 4073 7590 4085 7642
rect 4137 7590 8268 7642
rect 8320 7590 8332 7642
rect 8384 7590 8396 7642
rect 8448 7590 8460 7642
rect 8512 7590 8524 7642
rect 8576 7590 12707 7642
rect 12759 7590 12771 7642
rect 12823 7590 12835 7642
rect 12887 7590 12899 7642
rect 12951 7590 12963 7642
rect 13015 7590 17146 7642
rect 17198 7590 17210 7642
rect 17262 7590 17274 7642
rect 17326 7590 17338 7642
rect 17390 7590 17402 7642
rect 17454 7590 18860 7642
rect 1104 7568 18860 7590
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7377 7531 7435 7537
rect 7377 7528 7389 7531
rect 7156 7500 7389 7528
rect 7156 7488 7162 7500
rect 7377 7497 7389 7500
rect 7423 7497 7435 7531
rect 7377 7491 7435 7497
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 8662 7528 8668 7540
rect 8435 7500 8668 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 14090 7528 14096 7540
rect 12400 7500 14096 7528
rect 12400 7488 12406 7500
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 7558 7460 7564 7472
rect 3436 7432 7564 7460
rect 3436 7401 3464 7432
rect 7558 7420 7564 7432
rect 7616 7420 7622 7472
rect 12618 7460 12624 7472
rect 8588 7432 12624 7460
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7361 3479 7395
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 3421 7355 3479 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 5258 7392 5264 7404
rect 5219 7364 5264 7392
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6362 7392 6368 7404
rect 6043 7364 6368 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 8588 7401 8616 7432
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6696 7364 7205 7392
rect 6696 7352 6702 7364
rect 7193 7361 7205 7364
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7361 8631 7395
rect 9214 7392 9220 7404
rect 9175 7364 9220 7392
rect 8573 7355 8631 7361
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7392 10563 7395
rect 10686 7392 10692 7404
rect 10551 7364 10692 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11204 7364 11713 7392
rect 11204 7352 11210 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 12250 7352 12256 7404
rect 12308 7392 12314 7404
rect 14921 7395 14979 7401
rect 14921 7392 14933 7395
rect 12308 7364 14933 7392
rect 12308 7352 12314 7364
rect 14921 7361 14933 7364
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 6454 7324 6460 7336
rect 2179 7296 6460 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 9398 7324 9404 7336
rect 6779 7296 9404 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 11480 7296 12357 7324
rect 11480 7284 11486 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12345 7287 12403 7293
rect 12452 7296 13001 7324
rect 2777 7259 2835 7265
rect 2777 7225 2789 7259
rect 2823 7256 2835 7259
rect 7006 7256 7012 7268
rect 2823 7228 7012 7256
rect 2823 7225 2835 7228
rect 2777 7219 2835 7225
rect 7006 7216 7012 7228
rect 7064 7216 7070 7268
rect 11698 7216 11704 7268
rect 11756 7256 11762 7268
rect 12452 7256 12480 7296
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 17497 7327 17555 7333
rect 17497 7324 17509 7327
rect 13964 7296 17509 7324
rect 13964 7284 13970 7296
rect 17497 7293 17509 7296
rect 17543 7293 17555 7327
rect 17497 7287 17555 7293
rect 14277 7259 14335 7265
rect 14277 7256 14289 7259
rect 11756 7228 12480 7256
rect 12544 7228 14289 7256
rect 11756 7216 11762 7228
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 4212 7160 5825 7188
rect 4212 7148 4218 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 9309 7191 9367 7197
rect 9309 7157 9321 7191
rect 9355 7188 9367 7191
rect 9398 7188 9404 7200
rect 9355 7160 9404 7188
rect 9355 7157 9367 7160
rect 9309 7151 9367 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12544 7188 12572 7228
rect 14277 7225 14289 7228
rect 14323 7225 14335 7259
rect 14277 7219 14335 7225
rect 14918 7216 14924 7268
rect 14976 7256 14982 7268
rect 15565 7259 15623 7265
rect 15565 7256 15577 7259
rect 14976 7228 15577 7256
rect 14976 7216 14982 7228
rect 15565 7225 15577 7228
rect 15611 7225 15623 7259
rect 15565 7219 15623 7225
rect 16850 7188 16856 7200
rect 12124 7160 12572 7188
rect 16811 7160 16856 7188
rect 12124 7148 12130 7160
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 18138 7188 18144 7200
rect 18099 7160 18144 7188
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 7466 6984 7472 6996
rect 5215 6956 7472 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 9214 6984 9220 6996
rect 9175 6956 9220 6984
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 13320 6956 15577 6984
rect 13320 6944 13326 6956
rect 15565 6953 15577 6956
rect 15611 6953 15623 6987
rect 15565 6947 15623 6953
rect 7282 6916 7288 6928
rect 5736 6888 7288 6916
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6848 2191 6851
rect 4338 6848 4344 6860
rect 2179 6820 4344 6848
rect 2179 6817 2191 6820
rect 2133 6811 2191 6817
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 5534 6848 5540 6860
rect 4448 6820 5540 6848
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 4448 6780 4476 6820
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 3467 6752 4476 6780
rect 4525 6783 4583 6789
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 5736 6780 5764 6888
rect 7282 6876 7288 6888
rect 7340 6876 7346 6928
rect 16209 6919 16267 6925
rect 16209 6916 16221 6919
rect 14108 6888 16221 6916
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6848 6515 6851
rect 7837 6851 7895 6857
rect 6503 6820 7696 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 4571 6752 5764 6780
rect 5813 6783 5871 6789
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6914 6780 6920 6792
rect 5859 6752 6408 6780
rect 6875 6752 6920 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 2792 6644 2820 6743
rect 6178 6712 6184 6724
rect 3528 6684 6184 6712
rect 3528 6644 3556 6684
rect 6178 6672 6184 6684
rect 6236 6672 6242 6724
rect 6380 6712 6408 6752
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7668 6780 7696 6820
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 9490 6848 9496 6860
rect 7883 6820 9496 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10318 6848 10324 6860
rect 9907 6820 10324 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10505 6851 10563 6857
rect 10505 6817 10517 6851
rect 10551 6848 10563 6851
rect 10594 6848 10600 6860
rect 10551 6820 10600 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10928 6820 10977 6848
rect 10928 6808 10934 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11296 6820 11621 6848
rect 11296 6808 11302 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 11848 6820 12909 6848
rect 11848 6808 11854 6820
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 14108 6848 14136 6888
rect 16209 6885 16221 6888
rect 16255 6885 16267 6919
rect 16209 6879 16267 6885
rect 16758 6876 16764 6928
rect 16816 6916 16822 6928
rect 16853 6919 16911 6925
rect 16853 6916 16865 6919
rect 16816 6888 16865 6916
rect 16816 6876 16822 6888
rect 16853 6885 16865 6888
rect 16899 6885 16911 6919
rect 16853 6879 16911 6885
rect 13504 6820 14136 6848
rect 13504 6808 13510 6820
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 18138 6848 18144 6860
rect 14516 6820 18144 6848
rect 14516 6808 14522 6820
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 8573 6783 8631 6789
rect 7668 6752 8156 6780
rect 8018 6712 8024 6724
rect 6380 6684 8024 6712
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 8128 6712 8156 6752
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 9950 6780 9956 6792
rect 8619 6752 9956 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 11572 6752 12265 6780
rect 11572 6740 11578 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 12253 6743 12311 6749
rect 12406 6752 13553 6780
rect 8938 6712 8944 6724
rect 8128 6684 8944 6712
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 12406 6712 12434 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 14148 6752 14289 6780
rect 14148 6740 14154 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 14921 6783 14979 6789
rect 14921 6780 14933 6783
rect 14700 6752 14933 6780
rect 14700 6740 14706 6752
rect 14921 6749 14933 6752
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 11940 6684 12434 6712
rect 11940 6672 11946 6684
rect 14826 6672 14832 6724
rect 14884 6712 14890 6724
rect 17512 6712 17540 6743
rect 14884 6684 17540 6712
rect 14884 6672 14890 6684
rect 2792 6616 3556 6644
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 5442 6644 5448 6656
rect 3660 6616 5448 6644
rect 3660 6604 3666 6616
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6730 6644 6736 6656
rect 5592 6616 6736 6644
rect 5592 6604 5598 6616
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 7101 6647 7159 6653
rect 7101 6644 7113 6647
rect 6880 6616 7113 6644
rect 6880 6604 6886 6616
rect 7101 6613 7113 6616
rect 7147 6613 7159 6647
rect 7101 6607 7159 6613
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 8168 6616 8401 6644
rect 8168 6604 8174 6616
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 8389 6607 8447 6613
rect 14366 6604 14372 6656
rect 14424 6644 14430 6656
rect 16758 6644 16764 6656
rect 14424 6616 16764 6644
rect 14424 6604 14430 6616
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 1104 6554 18860 6576
rect 1104 6502 3829 6554
rect 3881 6502 3893 6554
rect 3945 6502 3957 6554
rect 4009 6502 4021 6554
rect 4073 6502 4085 6554
rect 4137 6502 8268 6554
rect 8320 6502 8332 6554
rect 8384 6502 8396 6554
rect 8448 6502 8460 6554
rect 8512 6502 8524 6554
rect 8576 6502 12707 6554
rect 12759 6502 12771 6554
rect 12823 6502 12835 6554
rect 12887 6502 12899 6554
rect 12951 6502 12963 6554
rect 13015 6502 17146 6554
rect 17198 6502 17210 6554
rect 17262 6502 17274 6554
rect 17326 6502 17338 6554
rect 17390 6502 17402 6554
rect 17454 6502 18860 6554
rect 1104 6480 18860 6502
rect 2746 6412 3832 6440
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 2746 6304 2774 6412
rect 2639 6276 2774 6304
rect 3804 6304 3832 6412
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 3936 6412 6040 6440
rect 3936 6400 3942 6412
rect 3970 6332 3976 6384
rect 4028 6372 4034 6384
rect 5902 6372 5908 6384
rect 4028 6344 5908 6372
rect 4028 6332 4034 6344
rect 5902 6332 5908 6344
rect 5960 6332 5966 6384
rect 6012 6372 6040 6412
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 12713 6443 12771 6449
rect 12713 6440 12725 6443
rect 12676 6412 12725 6440
rect 12676 6400 12682 6412
rect 12713 6409 12725 6412
rect 12759 6409 12771 6443
rect 12713 6403 12771 6409
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13136 6412 14872 6440
rect 13136 6400 13142 6412
rect 6546 6372 6552 6384
rect 6012 6344 6552 6372
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 8846 6372 8852 6384
rect 7024 6344 8852 6372
rect 4246 6304 4252 6316
rect 3804 6276 4252 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 6638 6304 6644 6316
rect 5307 6276 6644 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 7024 6313 7052 6344
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 12434 6332 12440 6384
rect 12492 6372 12498 6384
rect 12492 6344 14228 6372
rect 12492 6332 12498 6344
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7009 6267 7067 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 9582 6304 9588 6316
rect 8803 6276 9588 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 3878 6236 3884 6248
rect 3839 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4430 6196 4436 6248
rect 4488 6236 4494 6248
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4488 6208 4997 6236
rect 4488 6196 4494 6208
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 4985 6199 5043 6205
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7668 6236 7696 6267
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6304 10103 6307
rect 10134 6304 10140 6316
rect 10091 6276 10140 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10468 6276 10517 6304
rect 10468 6264 10474 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 10505 6267 10563 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11848 6276 11897 6304
rect 11848 6264 11854 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 13446 6304 13452 6316
rect 13407 6276 13452 6304
rect 11885 6267 11943 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 14200 6313 14228 6344
rect 14844 6313 14872 6412
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 15068 6276 16865 6304
rect 15068 6264 15074 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 11716 6236 11744 6264
rect 7340 6208 11744 6236
rect 7340 6196 7346 6208
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 13780 6208 13825 6236
rect 13780 6196 13786 6208
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 14516 6208 16129 6236
rect 14516 6196 14522 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6168 2007 6171
rect 5997 6171 6055 6177
rect 1995 6140 4660 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 3970 6100 3976 6112
rect 3283 6072 3976 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 4632 6100 4660 6140
rect 5997 6137 6009 6171
rect 6043 6168 6055 6171
rect 6914 6168 6920 6180
rect 6043 6140 6920 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 7837 6171 7895 6177
rect 7837 6137 7849 6171
rect 7883 6168 7895 6171
rect 8846 6168 8852 6180
rect 7883 6140 8852 6168
rect 7883 6137 7895 6140
rect 7837 6131 7895 6137
rect 8846 6128 8852 6140
rect 8904 6128 8910 6180
rect 9401 6171 9459 6177
rect 9401 6137 9413 6171
rect 9447 6168 9459 6171
rect 10042 6168 10048 6180
rect 9447 6140 10048 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 15473 6171 15531 6177
rect 15473 6168 15485 6171
rect 10152 6140 12020 6168
rect 5350 6100 5356 6112
rect 4632 6072 5356 6100
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 10152 6100 10180 6140
rect 11992 6112 12020 6140
rect 13648 6140 15485 6168
rect 13648 6112 13676 6140
rect 15473 6137 15485 6140
rect 15519 6137 15531 6171
rect 15473 6131 15531 6137
rect 7984 6072 10180 6100
rect 7984 6060 7990 6072
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 11572 6072 11897 6100
rect 11572 6060 11578 6072
rect 11885 6069 11897 6072
rect 11931 6069 11943 6103
rect 11885 6063 11943 6069
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 12032 6072 12173 6100
rect 12032 6060 12038 6072
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 12161 6063 12219 6069
rect 13630 6060 13636 6112
rect 13688 6060 13694 6112
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4764 5868 4813 5896
rect 4764 5856 4770 5868
rect 4801 5865 4813 5868
rect 4847 5865 4859 5899
rect 6638 5896 6644 5908
rect 4801 5859 4859 5865
rect 4908 5868 6224 5896
rect 6599 5868 6644 5896
rect 4522 5788 4528 5840
rect 4580 5828 4586 5840
rect 4908 5828 4936 5868
rect 4580 5800 4936 5828
rect 6196 5828 6224 5868
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 7745 5899 7803 5905
rect 7745 5865 7757 5899
rect 7791 5865 7803 5899
rect 7745 5859 7803 5865
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 9214 5896 9220 5908
rect 8619 5868 9220 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 7190 5828 7196 5840
rect 6196 5800 7196 5828
rect 4580 5788 4586 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 7377 5831 7435 5837
rect 7377 5828 7389 5831
rect 7340 5800 7389 5828
rect 7340 5788 7346 5800
rect 7377 5797 7389 5800
rect 7423 5797 7435 5831
rect 7377 5791 7435 5797
rect 1946 5720 1952 5772
rect 2004 5760 2010 5772
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 2004 5732 3341 5760
rect 2004 5720 2010 5732
rect 3329 5729 3341 5732
rect 3375 5760 3387 5763
rect 4338 5760 4344 5772
rect 3375 5732 4344 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 7760 5760 7788 5859
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 10597 5899 10655 5905
rect 10597 5896 10609 5899
rect 9916 5868 10609 5896
rect 9916 5856 9922 5868
rect 10597 5865 10609 5868
rect 10643 5865 10655 5899
rect 10597 5859 10655 5865
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 12584 5868 13553 5896
rect 12584 5856 12590 5868
rect 13541 5865 13553 5868
rect 13587 5865 13599 5899
rect 13541 5859 13599 5865
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 15565 5899 15623 5905
rect 15565 5896 15577 5899
rect 14792 5868 15577 5896
rect 14792 5856 14798 5868
rect 15565 5865 15577 5868
rect 15611 5865 15623 5899
rect 15565 5859 15623 5865
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 10137 5831 10195 5837
rect 10137 5828 10149 5831
rect 10008 5800 10149 5828
rect 10008 5788 10014 5800
rect 10137 5797 10149 5800
rect 10183 5797 10195 5831
rect 10137 5791 10195 5797
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 14921 5831 14979 5837
rect 14921 5828 14933 5831
rect 14056 5800 14933 5828
rect 14056 5788 14062 5800
rect 14921 5797 14933 5800
rect 14967 5797 14979 5831
rect 14921 5791 14979 5797
rect 6288 5732 7788 5760
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 2958 5652 2964 5704
rect 3016 5652 3022 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3752 5664 3985 5692
rect 3752 5652 3758 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 4982 5692 4988 5704
rect 4939 5664 4988 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5258 5692 5264 5704
rect 5215 5664 5264 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5626 5692 5632 5704
rect 5587 5664 5632 5692
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 6288 5692 6316 5732
rect 5951 5664 6316 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 1854 5624 1860 5636
rect 1815 5596 1860 5624
rect 1854 5584 1860 5596
rect 1912 5584 1918 5636
rect 5920 5624 5948 5655
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 9088 5664 9137 5692
rect 9088 5652 9094 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9398 5692 9404 5704
rect 9359 5664 9404 5692
rect 9125 5655 9183 5661
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 9968 5624 9996 5788
rect 11514 5760 11520 5772
rect 11475 5732 11520 5760
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 13412 5732 14289 5760
rect 13412 5720 13418 5732
rect 14277 5729 14289 5732
rect 14323 5729 14335 5763
rect 14277 5723 14335 5729
rect 11238 5692 11244 5704
rect 11199 5664 11244 5692
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 12618 5652 12624 5704
rect 12676 5652 12682 5704
rect 4172 5596 5948 5624
rect 6012 5596 9996 5624
rect 4172 5565 4200 5596
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5525 4215 5559
rect 4614 5556 4620 5568
rect 4575 5528 4620 5556
rect 4157 5519 4215 5525
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 5258 5556 5264 5568
rect 4764 5528 5264 5556
rect 4764 5516 4770 5528
rect 5258 5516 5264 5528
rect 5316 5556 5322 5568
rect 6012 5556 6040 5596
rect 5316 5528 6040 5556
rect 7745 5559 7803 5565
rect 5316 5516 5322 5528
rect 7745 5525 7757 5559
rect 7791 5556 7803 5559
rect 7834 5556 7840 5568
rect 7791 5528 7840 5556
rect 7791 5525 7803 5528
rect 7745 5519 7803 5525
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 7929 5559 7987 5565
rect 7929 5525 7941 5559
rect 7975 5556 7987 5559
rect 8938 5556 8944 5568
rect 7975 5528 8944 5556
rect 7975 5525 7987 5528
rect 7929 5519 7987 5525
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 11882 5516 11888 5568
rect 11940 5556 11946 5568
rect 12989 5559 13047 5565
rect 12989 5556 13001 5559
rect 11940 5528 13001 5556
rect 11940 5516 11946 5528
rect 12989 5525 13001 5528
rect 13035 5556 13047 5559
rect 13354 5556 13360 5568
rect 13035 5528 13360 5556
rect 13035 5525 13047 5528
rect 12989 5519 13047 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 1104 5466 18860 5488
rect 1104 5414 3829 5466
rect 3881 5414 3893 5466
rect 3945 5414 3957 5466
rect 4009 5414 4021 5466
rect 4073 5414 4085 5466
rect 4137 5414 8268 5466
rect 8320 5414 8332 5466
rect 8384 5414 8396 5466
rect 8448 5414 8460 5466
rect 8512 5414 8524 5466
rect 8576 5414 12707 5466
rect 12759 5414 12771 5466
rect 12823 5414 12835 5466
rect 12887 5414 12899 5466
rect 12951 5414 12963 5466
rect 13015 5414 17146 5466
rect 17198 5414 17210 5466
rect 17262 5414 17274 5466
rect 17326 5414 17338 5466
rect 17390 5414 17402 5466
rect 17454 5414 18860 5466
rect 1104 5392 18860 5414
rect 2746 5324 4292 5352
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 1946 5216 1952 5228
rect 1627 5188 1952 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2746 5148 2774 5324
rect 4264 5284 4292 5324
rect 5258 5312 5264 5364
rect 5316 5312 5322 5364
rect 5350 5312 5356 5364
rect 5408 5312 5414 5364
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 5626 5352 5632 5364
rect 5583 5324 5632 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 7524 5324 7757 5352
rect 7524 5312 7530 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 7745 5315 7803 5321
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11296 5324 12081 5352
rect 11296 5312 11302 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12069 5315 12127 5321
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12897 5355 12955 5361
rect 12299 5324 12434 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 4798 5284 4804 5296
rect 4264 5256 4804 5284
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 5276 5247 5304 5312
rect 5368 5247 5396 5312
rect 7374 5284 7380 5296
rect 6748 5256 7380 5284
rect 5261 5241 5319 5247
rect 4157 5228 4215 5231
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3697 5219 3755 5225
rect 3697 5216 3709 5219
rect 3660 5188 3709 5216
rect 3660 5176 3666 5188
rect 3697 5185 3709 5188
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 4154 5176 4160 5228
rect 4212 5222 4218 5228
rect 4212 5194 4251 5222
rect 4341 5219 4399 5225
rect 4212 5176 4218 5194
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 5151 5219 5209 5225
rect 5151 5216 5163 5219
rect 4341 5179 4399 5185
rect 5148 5185 5163 5216
rect 5197 5185 5209 5219
rect 5261 5207 5273 5241
rect 5307 5207 5319 5241
rect 5261 5201 5319 5207
rect 5353 5241 5411 5247
rect 5353 5207 5365 5241
rect 5399 5207 5411 5241
rect 6748 5225 6776 5256
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 7834 5284 7840 5296
rect 7484 5256 7840 5284
rect 5353 5201 5411 5207
rect 6733 5219 6791 5225
rect 5148 5179 5209 5185
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 7484 5216 7512 5256
rect 7834 5244 7840 5256
rect 7892 5244 7898 5296
rect 7331 5188 7512 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 2455 5120 2774 5148
rect 4356 5148 4384 5179
rect 4982 5148 4988 5160
rect 4356 5120 4988 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 4982 5108 4988 5120
rect 5040 5148 5046 5160
rect 5148 5148 5176 5179
rect 7300 5148 7328 5179
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 8665 5219 8723 5225
rect 7616 5188 7661 5216
rect 7616 5176 7622 5188
rect 8665 5185 8677 5219
rect 8711 5216 8723 5219
rect 8754 5216 8760 5228
rect 8711 5188 8760 5216
rect 8711 5185 8723 5188
rect 8665 5179 8723 5185
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9824 5188 9873 5216
rect 9824 5176 9830 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 11882 5216 11888 5228
rect 11747 5188 11888 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 12406 5216 12434 5324
rect 12897 5321 12909 5355
rect 12943 5352 12955 5355
rect 13446 5352 13452 5364
rect 12943 5324 13452 5352
rect 12943 5321 12955 5324
rect 12897 5315 12955 5321
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 12406 5188 12725 5216
rect 12713 5185 12725 5188
rect 12759 5185 12771 5219
rect 13354 5216 13360 5228
rect 13315 5188 13360 5216
rect 12713 5179 12771 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14550 5176 14556 5228
rect 14608 5216 14614 5228
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 14608 5188 14657 5216
rect 14608 5176 14614 5188
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 15252 5188 15301 5216
rect 15252 5176 15258 5188
rect 15289 5185 15301 5188
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 5040 5120 5212 5148
rect 5040 5108 5046 5120
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 5074 5080 5080 5092
rect 3099 5052 5080 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 5184 5080 5212 5120
rect 5368 5120 7328 5148
rect 5368 5080 5396 5120
rect 7374 5080 7380 5092
rect 5184 5052 5396 5080
rect 7335 5052 7380 5080
rect 7374 5040 7380 5052
rect 7432 5040 7438 5092
rect 7469 5083 7527 5089
rect 7469 5049 7481 5083
rect 7515 5080 7527 5083
rect 8018 5080 8024 5092
rect 7515 5052 8024 5080
rect 7515 5049 7527 5052
rect 7469 5043 7527 5049
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 4338 5012 4344 5024
rect 4299 4984 4344 5012
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 5902 5012 5908 5024
rect 4571 4984 5908 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 11756 4984 12081 5012
rect 11756 4972 11762 4984
rect 12069 4981 12081 4984
rect 12115 4981 12127 5015
rect 12069 4975 12127 4981
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 13541 5015 13599 5021
rect 13541 5012 13553 5015
rect 13412 4984 13553 5012
rect 13412 4972 13418 4984
rect 13541 4981 13553 4984
rect 13587 4981 13599 5015
rect 13541 4975 13599 4981
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 4172 4780 5641 4808
rect 4172 4749 4200 4780
rect 5629 4777 5641 4780
rect 5675 4808 5687 4811
rect 5902 4808 5908 4820
rect 5675 4780 5908 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 9398 4808 9404 4820
rect 9355 4780 9404 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12676 4780 12817 4808
rect 12676 4768 12682 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 12805 4771 12863 4777
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13722 4808 13728 4820
rect 13587 4780 13728 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 4157 4743 4215 4749
rect 4157 4709 4169 4743
rect 4203 4709 4215 4743
rect 4157 4703 4215 4709
rect 4985 4743 5043 4749
rect 4985 4709 4997 4743
rect 5031 4740 5043 4743
rect 6086 4740 6092 4752
rect 5031 4712 6092 4740
rect 5031 4709 5043 4712
rect 4985 4703 5043 4709
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 1673 4675 1731 4681
rect 1673 4672 1685 4675
rect 1636 4644 1685 4672
rect 1636 4632 1642 4644
rect 1673 4641 1685 4644
rect 1719 4672 1731 4675
rect 1719 4644 3648 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 3050 4564 3056 4616
rect 3108 4564 3114 4616
rect 3620 4604 3648 4644
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 5000 4672 5028 4703
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 9306 4672 9312 4684
rect 3752 4644 5028 4672
rect 6840 4644 9312 4672
rect 3752 4632 3758 4644
rect 6840 4613 6868 4644
rect 9306 4632 9312 4644
rect 9364 4672 9370 4684
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 9364 4644 10517 4672
rect 9364 4632 9370 4644
rect 10505 4641 10517 4644
rect 10551 4672 10563 4675
rect 11238 4672 11244 4684
rect 10551 4644 11244 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 3620 4576 6837 4604
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 8938 4564 8944 4616
rect 8996 4604 9002 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8996 4576 9137 4604
rect 8996 4564 9002 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9214 4564 9220 4616
rect 9272 4604 9278 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9272 4576 9873 4604
rect 9272 4564 9278 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12584 4576 12725 4604
rect 12584 4564 12590 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 12713 4567 12771 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 1946 4536 1952 4548
rect 1907 4508 1952 4536
rect 1946 4496 1952 4508
rect 2004 4496 2010 4548
rect 4433 4539 4491 4545
rect 4433 4536 4445 4539
rect 3436 4508 4445 4536
rect 3436 4477 3464 4508
rect 4433 4505 4445 4508
rect 4479 4536 4491 4539
rect 5350 4536 5356 4548
rect 4479 4508 5356 4536
rect 4479 4505 4491 4508
rect 4433 4499 4491 4505
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 5445 4539 5503 4545
rect 5445 4505 5457 4539
rect 5491 4536 5503 4539
rect 5534 4536 5540 4548
rect 5491 4508 5540 4536
rect 5491 4505 5503 4508
rect 5445 4499 5503 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 7098 4536 7104 4548
rect 7059 4508 7104 4536
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 8662 4536 8668 4548
rect 8326 4508 8668 4536
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 10781 4539 10839 4545
rect 10781 4505 10793 4539
rect 10827 4505 10839 4539
rect 10781 4499 10839 4505
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4437 3479 4471
rect 3421 4431 3479 4437
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 3568 4440 3985 4468
rect 3568 4428 3574 4440
rect 3973 4437 3985 4440
rect 4019 4437 4031 4471
rect 3973 4431 4031 4437
rect 5626 4428 5632 4480
rect 5684 4477 5690 4480
rect 5684 4471 5703 4477
rect 5691 4437 5703 4471
rect 5810 4468 5816 4480
rect 5771 4440 5816 4468
rect 5684 4431 5703 4437
rect 5684 4428 5690 4431
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8573 4471 8631 4477
rect 8573 4468 8585 4471
rect 8076 4440 8585 4468
rect 8076 4428 8082 4440
rect 8573 4437 8585 4440
rect 8619 4437 8631 4471
rect 8573 4431 8631 4437
rect 10045 4471 10103 4477
rect 10045 4437 10057 4471
rect 10091 4468 10103 4471
rect 10796 4468 10824 4499
rect 11790 4496 11796 4548
rect 11848 4496 11854 4548
rect 12250 4468 12256 4480
rect 10091 4440 10824 4468
rect 12211 4440 12256 4468
rect 10091 4437 10103 4440
rect 10045 4431 10103 4437
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 1104 4378 18860 4400
rect 1104 4326 3829 4378
rect 3881 4326 3893 4378
rect 3945 4326 3957 4378
rect 4009 4326 4021 4378
rect 4073 4326 4085 4378
rect 4137 4326 8268 4378
rect 8320 4326 8332 4378
rect 8384 4326 8396 4378
rect 8448 4326 8460 4378
rect 8512 4326 8524 4378
rect 8576 4326 12707 4378
rect 12759 4326 12771 4378
rect 12823 4326 12835 4378
rect 12887 4326 12899 4378
rect 12951 4326 12963 4378
rect 13015 4326 17146 4378
rect 17198 4326 17210 4378
rect 17262 4326 17274 4378
rect 17326 4326 17338 4378
rect 17390 4326 17402 4378
rect 17454 4326 18860 4378
rect 1104 4304 18860 4326
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 7466 4264 7472 4276
rect 5408 4236 7472 4264
rect 5408 4224 5414 4236
rect 7466 4224 7472 4236
rect 7524 4264 7530 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7524 4236 7573 4264
rect 7524 4224 7530 4236
rect 7561 4233 7573 4236
rect 7607 4264 7619 4267
rect 7607 4236 8156 4264
rect 7607 4233 7619 4236
rect 7561 4227 7619 4233
rect 5276 4168 7144 4196
rect 5276 4140 5304 4168
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 2501 4131 2559 4137
rect 2501 4128 2513 4131
rect 1820 4100 2513 4128
rect 1820 4088 1826 4100
rect 2501 4097 2513 4100
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 3016 4100 3065 4128
rect 3016 4088 3022 4100
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3602 4128 3608 4140
rect 3191 4100 3608 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 4614 4128 4620 4140
rect 3927 4100 4620 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5258 4128 5264 4140
rect 5215 4100 5264 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 5534 4128 5540 4140
rect 5408 4100 5453 4128
rect 5495 4100 5540 4128
rect 5408 4088 5414 4100
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6328 4100 6561 4128
rect 6328 4088 6334 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 7116 4060 7144 4168
rect 7374 4128 7380 4140
rect 7335 4100 7380 4128
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 8128 4137 8156 4236
rect 8389 4199 8447 4205
rect 8389 4165 8401 4199
rect 8435 4196 8447 4199
rect 12250 4196 12256 4208
rect 8435 4168 12256 4196
rect 8435 4165 8447 4168
rect 8389 4159 8447 4165
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 7668 4060 7696 4091
rect 8018 4060 8024 4072
rect 7116 4032 8024 4060
rect 8018 4020 8024 4032
rect 8076 4060 8082 4072
rect 8220 4060 8248 4091
rect 8076 4032 8248 4060
rect 8076 4020 8082 4032
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 2317 3995 2375 4001
rect 2317 3992 2329 3995
rect 1912 3964 2329 3992
rect 1912 3952 1918 3964
rect 2317 3961 2329 3964
rect 2363 3961 2375 3995
rect 2317 3955 2375 3961
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 4430 3992 4436 4004
rect 4111 3964 4436 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 4430 3952 4436 3964
rect 4488 3952 4494 4004
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 5166 3992 5172 4004
rect 4755 3964 5172 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 8404 3992 8432 4159
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 8846 4128 8852 4140
rect 8807 4100 8852 4128
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 11790 4128 11796 4140
rect 11751 4100 11796 4128
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 12526 4128 12532 4140
rect 11940 4100 12532 4128
rect 11940 4088 11946 4100
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 9030 3992 9036 4004
rect 7432 3964 8432 3992
rect 8991 3964 9036 3992
rect 7432 3952 7438 3964
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 7282 3924 7288 3936
rect 7239 3896 7288 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 2004 3692 2329 3720
rect 2004 3680 2010 3692
rect 2317 3689 2329 3692
rect 2363 3689 2375 3723
rect 3050 3720 3056 3732
rect 3011 3692 3056 3720
rect 2317 3683 2375 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4948 3692 4997 3720
rect 4948 3680 4954 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 4985 3683 5043 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6641 3723 6699 3729
rect 6641 3689 6653 3723
rect 6687 3720 6699 3723
rect 7098 3720 7104 3732
rect 6687 3692 7104 3720
rect 6687 3689 6699 3692
rect 6641 3683 6699 3689
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 8662 3720 8668 3732
rect 8527 3692 8668 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 7469 3655 7527 3661
rect 7469 3621 7481 3655
rect 7515 3652 7527 3655
rect 9214 3652 9220 3664
rect 7515 3624 9220 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 3510 3584 3516 3596
rect 2516 3556 3516 3584
rect 2516 3525 2544 3556
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 5736 3556 8616 3584
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3602 3516 3608 3528
rect 3191 3488 3608 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3602 3476 3608 3488
rect 3660 3516 3666 3528
rect 4154 3516 4160 3528
rect 3660 3488 4160 3516
rect 3660 3476 3666 3488
rect 4154 3476 4160 3488
rect 4212 3516 4218 3528
rect 5736 3516 5764 3556
rect 4212 3488 5764 3516
rect 4212 3476 4218 3488
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 8588 3525 8616 3556
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 5868 3488 6469 3516
rect 5868 3476 5874 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 11882 3516 11888 3528
rect 8619 3488 11888 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 7101 3451 7159 3457
rect 7101 3448 7113 3451
rect 5960 3420 7113 3448
rect 5960 3408 5966 3420
rect 7101 3417 7113 3420
rect 7147 3417 7159 3451
rect 7101 3411 7159 3417
rect 7317 3451 7375 3457
rect 7317 3417 7329 3451
rect 7363 3448 7375 3451
rect 8110 3448 8116 3460
rect 7363 3420 8116 3448
rect 7363 3417 7375 3420
rect 7317 3411 7375 3417
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 1104 3290 18860 3312
rect 1104 3238 3829 3290
rect 3881 3238 3893 3290
rect 3945 3238 3957 3290
rect 4009 3238 4021 3290
rect 4073 3238 4085 3290
rect 4137 3238 8268 3290
rect 8320 3238 8332 3290
rect 8384 3238 8396 3290
rect 8448 3238 8460 3290
rect 8512 3238 8524 3290
rect 8576 3238 12707 3290
rect 12759 3238 12771 3290
rect 12823 3238 12835 3290
rect 12887 3238 12899 3290
rect 12951 3238 12963 3290
rect 13015 3238 17146 3290
rect 17198 3238 17210 3290
rect 17262 3238 17274 3290
rect 17326 3238 17338 3290
rect 17390 3238 17402 3290
rect 17454 3238 18860 3290
rect 1104 3216 18860 3238
rect 5445 3179 5503 3185
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 5626 3176 5632 3188
rect 5491 3148 5632 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 5316 3012 5365 3040
rect 5316 3000 5322 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 5500 3012 5549 3040
rect 5500 3000 5506 3012
rect 5537 3009 5549 3012
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 1104 2202 18860 2224
rect 1104 2150 3829 2202
rect 3881 2150 3893 2202
rect 3945 2150 3957 2202
rect 4009 2150 4021 2202
rect 4073 2150 4085 2202
rect 4137 2150 8268 2202
rect 8320 2150 8332 2202
rect 8384 2150 8396 2202
rect 8448 2150 8460 2202
rect 8512 2150 8524 2202
rect 8576 2150 12707 2202
rect 12759 2150 12771 2202
rect 12823 2150 12835 2202
rect 12887 2150 12899 2202
rect 12951 2150 12963 2202
rect 13015 2150 17146 2202
rect 17198 2150 17210 2202
rect 17262 2150 17274 2202
rect 17326 2150 17338 2202
rect 17390 2150 17402 2202
rect 17454 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 12808 8236 12860 8288
rect 14924 8236 14976 8288
rect 5264 7964 5316 8016
rect 8668 7964 8720 8016
rect 8576 7896 8628 7948
rect 9220 7896 9272 7948
rect 7288 7760 7340 7812
rect 7656 7760 7708 7812
rect 4620 7692 4672 7744
rect 7932 7692 7984 7744
rect 8392 7692 8444 7744
rect 8852 7692 8904 7744
rect 12900 7692 12952 7744
rect 14648 7692 14700 7744
rect 3829 7590 3881 7642
rect 3893 7590 3945 7642
rect 3957 7590 4009 7642
rect 4021 7590 4073 7642
rect 4085 7590 4137 7642
rect 8268 7590 8320 7642
rect 8332 7590 8384 7642
rect 8396 7590 8448 7642
rect 8460 7590 8512 7642
rect 8524 7590 8576 7642
rect 12707 7590 12759 7642
rect 12771 7590 12823 7642
rect 12835 7590 12887 7642
rect 12899 7590 12951 7642
rect 12963 7590 13015 7642
rect 17146 7590 17198 7642
rect 17210 7590 17262 7642
rect 17274 7590 17326 7642
rect 17338 7590 17390 7642
rect 17402 7590 17454 7642
rect 7104 7488 7156 7540
rect 8668 7488 8720 7540
rect 12348 7488 12400 7540
rect 14096 7488 14148 7540
rect 7564 7420 7616 7472
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 6368 7352 6420 7404
rect 6644 7352 6696 7404
rect 12624 7420 12676 7472
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 10692 7352 10744 7404
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11152 7352 11204 7404
rect 12256 7352 12308 7404
rect 6460 7284 6512 7336
rect 9404 7284 9456 7336
rect 11428 7284 11480 7336
rect 7012 7216 7064 7268
rect 11704 7216 11756 7268
rect 13912 7284 13964 7336
rect 4160 7148 4212 7200
rect 9404 7148 9456 7200
rect 12072 7148 12124 7200
rect 14924 7216 14976 7268
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 18144 7191 18196 7200
rect 18144 7157 18153 7191
rect 18153 7157 18187 7191
rect 18187 7157 18196 7191
rect 18144 7148 18196 7157
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 7472 6944 7524 6996
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 13268 6944 13320 6996
rect 4344 6808 4396 6860
rect 5540 6808 5592 6860
rect 7288 6876 7340 6928
rect 6920 6783 6972 6792
rect 6184 6672 6236 6724
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 9496 6808 9548 6860
rect 10324 6808 10376 6860
rect 10600 6808 10652 6860
rect 10876 6808 10928 6860
rect 11244 6808 11296 6860
rect 11796 6808 11848 6860
rect 13452 6808 13504 6860
rect 16764 6876 16816 6928
rect 14464 6808 14516 6860
rect 18144 6808 18196 6860
rect 8024 6672 8076 6724
rect 9956 6740 10008 6792
rect 11520 6740 11572 6792
rect 8944 6672 8996 6724
rect 11888 6672 11940 6724
rect 14096 6740 14148 6792
rect 14648 6740 14700 6792
rect 14832 6672 14884 6724
rect 3608 6604 3660 6656
rect 5448 6604 5500 6656
rect 5540 6604 5592 6656
rect 6736 6604 6788 6656
rect 6828 6604 6880 6656
rect 8116 6604 8168 6656
rect 14372 6604 14424 6656
rect 16764 6604 16816 6656
rect 3829 6502 3881 6554
rect 3893 6502 3945 6554
rect 3957 6502 4009 6554
rect 4021 6502 4073 6554
rect 4085 6502 4137 6554
rect 8268 6502 8320 6554
rect 8332 6502 8384 6554
rect 8396 6502 8448 6554
rect 8460 6502 8512 6554
rect 8524 6502 8576 6554
rect 12707 6502 12759 6554
rect 12771 6502 12823 6554
rect 12835 6502 12887 6554
rect 12899 6502 12951 6554
rect 12963 6502 13015 6554
rect 17146 6502 17198 6554
rect 17210 6502 17262 6554
rect 17274 6502 17326 6554
rect 17338 6502 17390 6554
rect 17402 6502 17454 6554
rect 3884 6400 3936 6452
rect 3976 6332 4028 6384
rect 5908 6332 5960 6384
rect 12624 6400 12676 6452
rect 13084 6400 13136 6452
rect 6552 6332 6604 6384
rect 4252 6264 4304 6316
rect 6644 6264 6696 6316
rect 8852 6332 8904 6384
rect 12440 6332 12492 6384
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 4436 6196 4488 6248
rect 7288 6196 7340 6248
rect 9588 6264 9640 6316
rect 10140 6264 10192 6316
rect 10416 6264 10468 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11796 6264 11848 6316
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 15016 6264 15068 6316
rect 13728 6239 13780 6248
rect 13728 6205 13737 6239
rect 13737 6205 13771 6239
rect 13771 6205 13780 6239
rect 13728 6196 13780 6205
rect 14464 6196 14516 6248
rect 3976 6060 4028 6112
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 6920 6128 6972 6180
rect 8852 6128 8904 6180
rect 10048 6128 10100 6180
rect 5356 6060 5408 6112
rect 7932 6060 7984 6112
rect 11520 6060 11572 6112
rect 11980 6060 12032 6112
rect 13636 6060 13688 6112
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 4712 5856 4764 5908
rect 6644 5899 6696 5908
rect 4528 5788 4580 5840
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 7196 5788 7248 5840
rect 7288 5788 7340 5840
rect 1952 5720 2004 5772
rect 4344 5720 4396 5772
rect 9220 5856 9272 5908
rect 9864 5856 9916 5908
rect 12532 5856 12584 5908
rect 14740 5856 14792 5908
rect 9956 5788 10008 5840
rect 14004 5788 14056 5840
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 2964 5652 3016 5704
rect 3700 5652 3752 5704
rect 4988 5652 5040 5704
rect 5264 5652 5316 5704
rect 5632 5695 5684 5704
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 1860 5627 1912 5636
rect 1860 5593 1869 5627
rect 1869 5593 1903 5627
rect 1903 5593 1912 5627
rect 1860 5584 1912 5593
rect 9036 5652 9088 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 13360 5720 13412 5772
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 12624 5652 12676 5704
rect 4620 5559 4672 5568
rect 4620 5525 4629 5559
rect 4629 5525 4663 5559
rect 4663 5525 4672 5559
rect 4620 5516 4672 5525
rect 4712 5516 4764 5568
rect 5264 5516 5316 5568
rect 7840 5516 7892 5568
rect 8944 5516 8996 5568
rect 11888 5516 11940 5568
rect 13360 5516 13412 5568
rect 3829 5414 3881 5466
rect 3893 5414 3945 5466
rect 3957 5414 4009 5466
rect 4021 5414 4073 5466
rect 4085 5414 4137 5466
rect 8268 5414 8320 5466
rect 8332 5414 8384 5466
rect 8396 5414 8448 5466
rect 8460 5414 8512 5466
rect 8524 5414 8576 5466
rect 12707 5414 12759 5466
rect 12771 5414 12823 5466
rect 12835 5414 12887 5466
rect 12899 5414 12951 5466
rect 12963 5414 13015 5466
rect 17146 5414 17198 5466
rect 17210 5414 17262 5466
rect 17274 5414 17326 5466
rect 17338 5414 17390 5466
rect 17402 5414 17454 5466
rect 1952 5176 2004 5228
rect 5264 5312 5316 5364
rect 5356 5312 5408 5364
rect 5632 5312 5684 5364
rect 7472 5312 7524 5364
rect 11244 5312 11296 5364
rect 4804 5244 4856 5296
rect 3608 5176 3660 5228
rect 4160 5225 4212 5228
rect 4160 5191 4169 5225
rect 4169 5191 4203 5225
rect 4203 5191 4212 5225
rect 4160 5176 4212 5191
rect 7380 5244 7432 5296
rect 7840 5244 7892 5296
rect 4988 5108 5040 5160
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 8760 5176 8812 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 9772 5176 9824 5228
rect 11888 5176 11940 5228
rect 13452 5312 13504 5364
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 14556 5176 14608 5228
rect 15200 5176 15252 5228
rect 5080 5040 5132 5092
rect 7380 5083 7432 5092
rect 7380 5049 7389 5083
rect 7389 5049 7423 5083
rect 7423 5049 7432 5083
rect 7380 5040 7432 5049
rect 8024 5040 8076 5092
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 4344 5015 4396 5024
rect 4344 4981 4353 5015
rect 4353 4981 4387 5015
rect 4387 4981 4396 5015
rect 4344 4972 4396 4981
rect 5908 4972 5960 5024
rect 11704 4972 11756 5024
rect 13360 4972 13412 5024
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 5908 4768 5960 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 9404 4768 9456 4820
rect 12624 4768 12676 4820
rect 13728 4768 13780 4820
rect 1584 4632 1636 4684
rect 3056 4564 3108 4616
rect 3700 4632 3752 4684
rect 6092 4700 6144 4752
rect 9312 4632 9364 4684
rect 11244 4632 11296 4684
rect 8944 4564 8996 4616
rect 9220 4564 9272 4616
rect 12532 4564 12584 4616
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 1952 4539 2004 4548
rect 1952 4505 1961 4539
rect 1961 4505 1995 4539
rect 1995 4505 2004 4539
rect 1952 4496 2004 4505
rect 5356 4496 5408 4548
rect 5540 4496 5592 4548
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 8668 4496 8720 4548
rect 3516 4428 3568 4480
rect 5632 4471 5684 4480
rect 5632 4437 5657 4471
rect 5657 4437 5684 4471
rect 5816 4471 5868 4480
rect 5632 4428 5684 4437
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 8024 4428 8076 4480
rect 11796 4496 11848 4548
rect 12256 4471 12308 4480
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 12256 4428 12308 4437
rect 3829 4326 3881 4378
rect 3893 4326 3945 4378
rect 3957 4326 4009 4378
rect 4021 4326 4073 4378
rect 4085 4326 4137 4378
rect 8268 4326 8320 4378
rect 8332 4326 8384 4378
rect 8396 4326 8448 4378
rect 8460 4326 8512 4378
rect 8524 4326 8576 4378
rect 12707 4326 12759 4378
rect 12771 4326 12823 4378
rect 12835 4326 12887 4378
rect 12899 4326 12951 4378
rect 12963 4326 13015 4378
rect 17146 4326 17198 4378
rect 17210 4326 17262 4378
rect 17274 4326 17326 4378
rect 17338 4326 17390 4378
rect 17402 4326 17454 4378
rect 5356 4224 5408 4276
rect 7472 4224 7524 4276
rect 1768 4088 1820 4140
rect 2964 4088 3016 4140
rect 3608 4088 3660 4140
rect 4620 4088 4672 4140
rect 5264 4088 5316 4140
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5540 4131 5592 4140
rect 5356 4088 5408 4097
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5540 4088 5592 4097
rect 6276 4088 6328 4140
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 8024 4020 8076 4072
rect 1860 3952 1912 4004
rect 4436 3952 4488 4004
rect 5172 3952 5224 4004
rect 7380 3952 7432 4004
rect 12256 4156 12308 4208
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12532 4088 12584 4140
rect 9036 3995 9088 4004
rect 9036 3961 9045 3995
rect 9045 3961 9079 3995
rect 9079 3961 9088 3995
rect 9036 3952 9088 3961
rect 7288 3884 7340 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 1952 3680 2004 3732
rect 3056 3723 3108 3732
rect 3056 3689 3065 3723
rect 3065 3689 3099 3723
rect 3099 3689 3108 3723
rect 3056 3680 3108 3689
rect 4896 3680 4948 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 7104 3680 7156 3732
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 8668 3680 8720 3732
rect 9220 3612 9272 3664
rect 3516 3544 3568 3596
rect 3608 3476 3660 3528
rect 4160 3476 4212 3528
rect 5816 3476 5868 3528
rect 11888 3476 11940 3528
rect 5908 3408 5960 3460
rect 8116 3408 8168 3460
rect 3829 3238 3881 3290
rect 3893 3238 3945 3290
rect 3957 3238 4009 3290
rect 4021 3238 4073 3290
rect 4085 3238 4137 3290
rect 8268 3238 8320 3290
rect 8332 3238 8384 3290
rect 8396 3238 8448 3290
rect 8460 3238 8512 3290
rect 8524 3238 8576 3290
rect 12707 3238 12759 3290
rect 12771 3238 12823 3290
rect 12835 3238 12887 3290
rect 12899 3238 12951 3290
rect 12963 3238 13015 3290
rect 17146 3238 17198 3290
rect 17210 3238 17262 3290
rect 17274 3238 17326 3290
rect 17338 3238 17390 3290
rect 17402 3238 17454 3290
rect 5632 3136 5684 3188
rect 5264 3000 5316 3052
rect 5448 3000 5500 3052
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 3829 2150 3881 2202
rect 3893 2150 3945 2202
rect 3957 2150 4009 2202
rect 4021 2150 4073 2202
rect 4085 2150 4137 2202
rect 8268 2150 8320 2202
rect 8332 2150 8384 2202
rect 8396 2150 8448 2202
rect 8460 2150 8512 2202
rect 8524 2150 8576 2202
rect 12707 2150 12759 2202
rect 12771 2150 12823 2202
rect 12835 2150 12887 2202
rect 12899 2150 12951 2202
rect 12963 2150 13015 2202
rect 17146 2150 17198 2202
rect 17210 2150 17262 2202
rect 17274 2150 17326 2202
rect 17338 2150 17390 2202
rect 17402 2150 17454 2202
<< metal2 >>
rect 4710 9200 4766 10000
rect 4802 9200 4858 10000
rect 4894 9200 4950 10000
rect 4986 9200 5042 10000
rect 5078 9200 5134 10000
rect 5170 9200 5226 10000
rect 5262 9200 5318 10000
rect 5354 9200 5410 10000
rect 5446 9200 5502 10000
rect 5538 9200 5594 10000
rect 5630 9200 5686 10000
rect 5722 9200 5778 10000
rect 5814 9200 5870 10000
rect 5906 9200 5962 10000
rect 5998 9200 6054 10000
rect 6090 9200 6146 10000
rect 6182 9200 6238 10000
rect 6274 9200 6330 10000
rect 6366 9200 6422 10000
rect 6458 9200 6514 10000
rect 6550 9200 6606 10000
rect 6642 9200 6698 10000
rect 6734 9200 6790 10000
rect 6826 9200 6882 10000
rect 6918 9200 6974 10000
rect 7010 9200 7066 10000
rect 7102 9200 7158 10000
rect 7194 9200 7250 10000
rect 7286 9200 7342 10000
rect 7378 9200 7434 10000
rect 7470 9200 7526 10000
rect 7562 9200 7618 10000
rect 7654 9200 7710 10000
rect 7746 9200 7802 10000
rect 7838 9200 7894 10000
rect 7930 9200 7986 10000
rect 8022 9200 8078 10000
rect 8114 9200 8170 10000
rect 8206 9200 8262 10000
rect 8298 9200 8354 10000
rect 8390 9200 8446 10000
rect 8482 9200 8538 10000
rect 8574 9200 8630 10000
rect 8666 9200 8722 10000
rect 8758 9200 8814 10000
rect 8850 9200 8906 10000
rect 8942 9200 8998 10000
rect 9034 9200 9090 10000
rect 9126 9200 9182 10000
rect 9218 9200 9274 10000
rect 9310 9200 9366 10000
rect 9402 9200 9458 10000
rect 9494 9200 9550 10000
rect 9586 9200 9642 10000
rect 9678 9200 9734 10000
rect 9770 9200 9826 10000
rect 9862 9200 9918 10000
rect 9954 9200 10010 10000
rect 10046 9200 10102 10000
rect 10138 9200 10194 10000
rect 10230 9200 10286 10000
rect 10322 9200 10378 10000
rect 10414 9200 10470 10000
rect 10506 9200 10562 10000
rect 10598 9200 10654 10000
rect 10690 9200 10746 10000
rect 10782 9200 10838 10000
rect 10874 9200 10930 10000
rect 10966 9200 11022 10000
rect 11058 9200 11114 10000
rect 11150 9200 11206 10000
rect 11242 9200 11298 10000
rect 11334 9200 11390 10000
rect 11426 9200 11482 10000
rect 11518 9200 11574 10000
rect 11610 9200 11666 10000
rect 11702 9200 11758 10000
rect 11794 9200 11850 10000
rect 11886 9200 11942 10000
rect 11978 9200 12034 10000
rect 12070 9200 12126 10000
rect 12162 9200 12218 10000
rect 12254 9200 12310 10000
rect 12346 9200 12402 10000
rect 12438 9200 12494 10000
rect 12530 9200 12586 10000
rect 12622 9200 12678 10000
rect 12714 9200 12770 10000
rect 12806 9200 12862 10000
rect 12898 9200 12954 10000
rect 12990 9200 13046 10000
rect 13082 9200 13138 10000
rect 13174 9200 13230 10000
rect 13266 9200 13322 10000
rect 13358 9200 13414 10000
rect 13450 9200 13506 10000
rect 13542 9200 13598 10000
rect 13634 9200 13690 10000
rect 13726 9200 13782 10000
rect 13818 9200 13874 10000
rect 13910 9200 13966 10000
rect 14002 9200 14058 10000
rect 14094 9200 14150 10000
rect 14186 9200 14242 10000
rect 14278 9200 14334 10000
rect 14370 9200 14426 10000
rect 14462 9200 14518 10000
rect 14554 9200 14610 10000
rect 14646 9200 14702 10000
rect 14738 9200 14794 10000
rect 14830 9200 14886 10000
rect 14922 9200 14978 10000
rect 15014 9200 15070 10000
rect 15106 9200 15162 10000
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 3829 7644 4137 7653
rect 3829 7642 3835 7644
rect 3891 7642 3915 7644
rect 3971 7642 3995 7644
rect 4051 7642 4075 7644
rect 4131 7642 4137 7644
rect 3891 7590 3893 7642
rect 4073 7590 4075 7642
rect 3829 7588 3835 7590
rect 3891 7588 3915 7590
rect 3971 7588 3995 7590
rect 4051 7588 4075 7590
rect 4131 7588 4137 7590
rect 3829 7579 4137 7588
rect 4632 7410 4660 7686
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 4690 1624 5646
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1780 4146 1808 4966
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1872 4010 1900 5578
rect 1964 5234 1992 5714
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1964 3738 1992 4490
rect 2976 4146 3004 5646
rect 3620 5234 3648 6598
rect 3829 6556 4137 6565
rect 3829 6554 3835 6556
rect 3891 6554 3915 6556
rect 3971 6554 3995 6556
rect 4051 6554 4075 6556
rect 4131 6554 4137 6556
rect 3891 6502 3893 6554
rect 4073 6502 4075 6554
rect 3829 6500 3835 6502
rect 3891 6500 3915 6502
rect 3971 6500 3995 6502
rect 4051 6500 4075 6502
rect 4131 6500 4137 6502
rect 3829 6491 4137 6500
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3896 6254 3924 6394
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3988 6118 4016 6326
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3712 4690 3740 5646
rect 3829 5468 4137 5477
rect 3829 5466 3835 5468
rect 3891 5466 3915 5468
rect 3971 5466 3995 5468
rect 4051 5466 4075 5468
rect 4131 5466 4137 5468
rect 3891 5414 3893 5466
rect 4073 5414 4075 5466
rect 3829 5412 3835 5414
rect 3891 5412 3915 5414
rect 3971 5412 3995 5414
rect 4051 5412 4075 5414
rect 4131 5412 4137 5414
rect 3829 5403 4137 5412
rect 4172 5234 4200 7142
rect 4342 6896 4398 6905
rect 4342 6831 4344 6840
rect 4396 6831 4398 6840
rect 4344 6802 4396 6808
rect 4250 6624 4306 6633
rect 4250 6559 4306 6568
rect 4264 6322 4292 6559
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4342 5808 4398 5817
rect 4342 5743 4344 5752
rect 4396 5743 4398 5752
rect 4344 5714 4396 5720
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3068 3738 3096 4558
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3528 3602 3556 4422
rect 3829 4380 4137 4389
rect 3829 4378 3835 4380
rect 3891 4378 3915 4380
rect 3971 4378 3995 4380
rect 4051 4378 4075 4380
rect 4131 4378 4137 4380
rect 3891 4326 3893 4378
rect 4073 4326 4075 4378
rect 3829 4324 3835 4326
rect 3891 4324 3915 4326
rect 3971 4324 3995 4326
rect 4051 4324 4075 4326
rect 4131 4324 4137 4326
rect 3829 4315 4137 4324
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3620 3534 3648 4082
rect 4172 3534 4200 5170
rect 4356 5030 4384 5714
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4448 4010 4476 6190
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5846 4568 6054
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4724 5574 4752 5850
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4632 4146 4660 5510
rect 4816 5302 4844 9200
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4908 3738 4936 9200
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5166 5028 5646
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5092 5098 5120 9200
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5184 4010 5212 9200
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5276 7410 5304 7958
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5368 6118 5396 9200
rect 5460 6662 5488 9200
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6662 5580 6802
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5644 6440 5672 9200
rect 5736 6633 5764 9200
rect 5920 6905 5948 9200
rect 5906 6896 5962 6905
rect 5906 6831 5962 6840
rect 5722 6624 5778 6633
rect 5722 6559 5778 6568
rect 5644 6412 5764 6440
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5262 5808 5318 5817
rect 5262 5743 5318 5752
rect 5276 5710 5304 5743
rect 5264 5704 5316 5710
rect 5632 5704 5684 5710
rect 5316 5664 5396 5692
rect 5264 5646 5316 5652
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5276 5370 5304 5510
rect 5368 5370 5396 5664
rect 5632 5646 5684 5652
rect 5644 5370 5672 5646
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5368 4282 5396 4490
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5368 4146 5396 4218
rect 5552 4146 5580 4490
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3829 3292 4137 3301
rect 3829 3290 3835 3292
rect 3891 3290 3915 3292
rect 3971 3290 3995 3292
rect 4051 3290 4075 3292
rect 4131 3290 4137 3292
rect 3891 3238 3893 3290
rect 4073 3238 4075 3290
rect 3829 3236 3835 3238
rect 3891 3236 3915 3238
rect 3971 3236 3995 3238
rect 4051 3236 4075 3238
rect 4131 3236 4137 3238
rect 3829 3227 4137 3236
rect 5276 3058 5304 4082
rect 5264 3052 5316 3058
rect 5368 3040 5396 4082
rect 5644 3194 5672 4422
rect 5736 3738 5764 6412
rect 5908 6384 5960 6390
rect 6012 6372 6040 9200
rect 5960 6344 6040 6372
rect 5908 6326 5960 6332
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4826 5948 4966
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5828 3534 5856 4422
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5920 3466 5948 4762
rect 6104 4758 6132 9200
rect 6196 6730 6224 9200
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6288 4146 6316 9200
rect 6380 7410 6408 9200
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6380 4826 6408 7346
rect 6472 7342 6500 9200
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6564 6390 6592 9200
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6656 6322 6684 7346
rect 6748 6662 6776 9200
rect 6840 6662 6868 9200
rect 7024 7274 7052 9200
rect 7116 7546 7144 9200
rect 7300 7970 7328 9200
rect 7208 7942 7328 7970
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 5914 6684 6258
rect 6932 6186 6960 6734
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 7208 5846 7236 7942
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7300 6934 7328 7754
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7300 5846 7328 6190
rect 7196 5840 7248 5846
rect 7288 5840 7340 5846
rect 7196 5782 7248 5788
rect 7286 5808 7288 5817
rect 7340 5808 7342 5817
rect 7286 5743 7342 5752
rect 7392 5302 7420 9200
rect 7576 7478 7604 9200
rect 7668 7818 7696 9200
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7852 7562 7880 9200
rect 7944 7750 7972 9200
rect 8128 7970 8156 9200
rect 8036 7942 8156 7970
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7668 7534 7880 7562
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7668 7290 7696 7534
rect 7484 7262 7696 7290
rect 7484 7002 7512 7262
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 8036 6730 8064 7942
rect 8220 7834 8248 9200
rect 8128 7806 8248 7834
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8128 6662 8156 7806
rect 8404 7750 8432 9200
rect 8496 7834 8524 9200
rect 8588 7954 8616 9200
rect 8680 8022 8708 9200
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8496 7806 8708 7834
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8268 7644 8576 7653
rect 8268 7642 8274 7644
rect 8330 7642 8354 7644
rect 8410 7642 8434 7644
rect 8490 7642 8514 7644
rect 8570 7642 8576 7644
rect 8330 7590 8332 7642
rect 8512 7590 8514 7642
rect 8268 7588 8274 7590
rect 8330 7588 8354 7590
rect 8410 7588 8434 7590
rect 8490 7588 8514 7590
rect 8570 7588 8576 7590
rect 8268 7579 8576 7588
rect 8680 7546 8708 7806
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8268 6556 8576 6565
rect 8268 6554 8274 6556
rect 8330 6554 8354 6556
rect 8410 6554 8434 6556
rect 8490 6554 8514 6556
rect 8570 6554 8576 6556
rect 8330 6502 8332 6554
rect 8512 6502 8514 6554
rect 8268 6500 8274 6502
rect 8330 6500 8354 6502
rect 8410 6500 8434 6502
rect 8490 6500 8514 6502
rect 8570 6500 8576 6502
rect 8268 6491 8576 6500
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7484 5370 7512 6258
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 7840 5568 7892 5574
rect 7944 5556 7972 6054
rect 7892 5528 7972 5556
rect 7840 5510 7892 5516
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7852 5302 7880 5510
rect 8268 5468 8576 5477
rect 8268 5466 8274 5468
rect 8330 5466 8354 5468
rect 8410 5466 8434 5468
rect 8490 5466 8514 5468
rect 8570 5466 8576 5468
rect 8330 5414 8332 5466
rect 8512 5414 8514 5466
rect 8268 5412 8274 5414
rect 8330 5412 8354 5414
rect 8410 5412 8434 5414
rect 8490 5412 8514 5414
rect 8570 5412 8576 5414
rect 8268 5403 8576 5412
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 8772 5234 8800 9200
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8864 6390 8892 7686
rect 8956 6730 8984 9200
rect 9048 7154 9076 9200
rect 9232 8106 9260 9200
rect 9324 8242 9352 9200
rect 9324 8214 9444 8242
rect 9232 8078 9352 8106
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9232 7410 9260 7890
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9048 7126 9168 7154
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 7564 5228 7616 5234
rect 7484 5188 7564 5216
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 7116 3738 7144 4490
rect 7392 4146 7420 5034
rect 7484 4282 7512 5188
rect 7564 5170 7616 5176
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 8036 4486 8064 5034
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7392 4010 7420 4082
rect 8036 4078 8064 4422
rect 8268 4380 8576 4389
rect 8268 4378 8274 4380
rect 8330 4378 8354 4380
rect 8410 4378 8434 4380
rect 8490 4378 8514 4380
rect 8570 4378 8576 4380
rect 8330 4326 8332 4378
rect 8512 4326 8514 4378
rect 8268 4324 8274 4326
rect 8330 4324 8354 4326
rect 8410 4324 8434 4326
rect 8490 4324 8514 4326
rect 8570 4324 8576 4326
rect 8268 4315 8576 4324
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7300 3738 7328 3878
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 8128 3466 8156 3878
rect 8680 3738 8708 4490
rect 8864 4146 8892 6122
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 4622 8984 5510
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 9048 4010 9076 5646
rect 9140 5234 9168 7126
rect 9232 7002 9260 7346
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9220 5908 9272 5914
rect 9324 5896 9352 8078
rect 9416 7342 9444 8214
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9272 5868 9352 5896
rect 9220 5850 9272 5856
rect 9416 5794 9444 7142
rect 9508 6866 9536 9200
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9600 6322 9628 9200
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9324 5766 9444 5794
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9324 4690 9352 5766
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 4826 9444 5646
rect 9784 5234 9812 9200
rect 9876 5914 9904 9200
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9968 5846 9996 6734
rect 10060 6186 10088 9200
rect 10152 6322 10180 9200
rect 10336 6866 10364 9200
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10428 6322 10456 9200
rect 10612 6866 10640 9200
rect 10704 7410 10732 9200
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10888 6866 10916 9200
rect 10980 7410 11008 9200
rect 11164 7410 11192 9200
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11256 6866 11284 9200
rect 11440 7342 11468 9200
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11532 6798 11560 9200
rect 11716 7274 11744 9200
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11808 6866 11836 9200
rect 11992 7154 12020 9200
rect 12084 7206 12112 9200
rect 12268 7410 12296 9200
rect 12360 7546 12388 9200
rect 12544 7698 12572 9200
rect 12452 7670 12572 7698
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 11900 7126 12020 7154
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11900 6730 11928 7126
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 12452 6390 12480 7670
rect 12636 7562 12664 9200
rect 12820 8294 12848 9200
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12912 7750 12940 9200
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12707 7644 13015 7653
rect 12707 7642 12713 7644
rect 12769 7642 12793 7644
rect 12849 7642 12873 7644
rect 12929 7642 12953 7644
rect 13009 7642 13015 7644
rect 12769 7590 12771 7642
rect 12951 7590 12953 7642
rect 12707 7588 12713 7590
rect 12769 7588 12793 7590
rect 12849 7588 12873 7590
rect 12929 7588 12953 7590
rect 13009 7588 13015 7590
rect 12707 7579 13015 7588
rect 12544 7534 12664 7562
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 11532 5778 11560 6054
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11256 5370 11284 5646
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 11256 4690 11284 5306
rect 11716 5030 11744 6258
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11808 4808 11836 6258
rect 11980 6112 12032 6118
rect 11900 6060 11980 6066
rect 11900 6054 12032 6060
rect 11900 6038 12020 6054
rect 11900 5574 11928 6038
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 12544 5914 12572 7534
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12636 6458 12664 7414
rect 12707 6556 13015 6565
rect 12707 6554 12713 6556
rect 12769 6554 12793 6556
rect 12849 6554 12873 6556
rect 12929 6554 12953 6556
rect 13009 6554 13015 6556
rect 12769 6502 12771 6554
rect 12951 6502 12953 6554
rect 12707 6500 12713 6502
rect 12769 6500 12793 6502
rect 12849 6500 12873 6502
rect 12929 6500 12953 6502
rect 13009 6500 13015 6502
rect 12707 6491 13015 6500
rect 13096 6458 13124 9200
rect 13188 7834 13216 9200
rect 13188 7806 13308 7834
rect 13280 7002 13308 7806
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 13372 5778 13400 9200
rect 13464 6866 13492 9200
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5234 11928 5510
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 12636 4826 12664 5646
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 12707 5468 13015 5477
rect 12707 5466 12713 5468
rect 12769 5466 12793 5468
rect 12849 5466 12873 5468
rect 12929 5466 12953 5468
rect 13009 5466 13015 5468
rect 12769 5414 12771 5466
rect 12951 5414 12953 5466
rect 12707 5412 12713 5414
rect 12769 5412 12793 5414
rect 12849 5412 12873 5414
rect 12929 5412 12953 5414
rect 13009 5412 13015 5414
rect 12707 5403 13015 5412
rect 13372 5234 13400 5510
rect 13464 5370 13492 6258
rect 13648 6118 13676 9200
rect 13740 6905 13768 9200
rect 13924 7342 13952 9200
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13726 6896 13782 6905
rect 13726 6831 13782 6840
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 12624 4820 12676 4826
rect 11808 4780 11928 4808
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 9232 3670 9260 4558
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11808 4146 11836 4490
rect 11900 4146 11928 4780
rect 12624 4762 12676 4768
rect 13372 4622 13400 4966
rect 13740 4826 13768 6190
rect 14016 5846 14044 9200
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14108 6798 14136 7482
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14200 6644 14228 9200
rect 14292 6746 14320 9200
rect 14476 6866 14504 9200
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14292 6718 14504 6746
rect 14372 6656 14424 6662
rect 14200 6616 14372 6644
rect 14372 6598 14424 6604
rect 14476 6254 14504 6718
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14568 5234 14596 9200
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 6798 14688 7686
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14752 5914 14780 9200
rect 14844 6730 14872 9200
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14936 7274 14964 8230
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 15028 6322 15056 9200
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 15120 5658 15148 9200
rect 17146 7644 17454 7653
rect 17146 7642 17152 7644
rect 17208 7642 17232 7644
rect 17288 7642 17312 7644
rect 17368 7642 17392 7644
rect 17448 7642 17454 7644
rect 17208 7590 17210 7642
rect 17390 7590 17392 7642
rect 17146 7588 17152 7590
rect 17208 7588 17232 7590
rect 17288 7588 17312 7590
rect 17368 7588 17392 7590
rect 17448 7588 17454 7590
rect 17146 7579 17454 7588
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 16764 6928 16816 6934
rect 16868 6905 16896 7142
rect 16764 6870 16816 6876
rect 16854 6896 16910 6905
rect 16776 6662 16804 6870
rect 18156 6866 18184 7142
rect 16854 6831 16910 6840
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 17146 6556 17454 6565
rect 17146 6554 17152 6556
rect 17208 6554 17232 6556
rect 17288 6554 17312 6556
rect 17368 6554 17392 6556
rect 17448 6554 17454 6556
rect 17208 6502 17210 6554
rect 17390 6502 17392 6554
rect 17146 6500 17152 6502
rect 17208 6500 17232 6502
rect 17288 6500 17312 6502
rect 17368 6500 17392 6502
rect 17448 6500 17454 6502
rect 17146 6491 17454 6500
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 15120 5630 15240 5658
rect 15212 5234 15240 5630
rect 17146 5468 17454 5477
rect 17146 5466 17152 5468
rect 17208 5466 17232 5468
rect 17288 5466 17312 5468
rect 17368 5466 17392 5468
rect 17448 5466 17454 5468
rect 17208 5414 17210 5466
rect 17390 5414 17392 5466
rect 17146 5412 17152 5414
rect 17208 5412 17232 5414
rect 17288 5412 17312 5414
rect 17368 5412 17392 5414
rect 17448 5412 17454 5414
rect 17146 5403 17454 5412
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12268 4214 12296 4422
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12544 4146 12572 4558
rect 12707 4380 13015 4389
rect 12707 4378 12713 4380
rect 12769 4378 12793 4380
rect 12849 4378 12873 4380
rect 12929 4378 12953 4380
rect 13009 4378 13015 4380
rect 12769 4326 12771 4378
rect 12951 4326 12953 4378
rect 12707 4324 12713 4326
rect 12769 4324 12793 4326
rect 12849 4324 12873 4326
rect 12929 4324 12953 4326
rect 13009 4324 13015 4326
rect 12707 4315 13015 4324
rect 17146 4380 17454 4389
rect 17146 4378 17152 4380
rect 17208 4378 17232 4380
rect 17288 4378 17312 4380
rect 17368 4378 17392 4380
rect 17448 4378 17454 4380
rect 17208 4326 17210 4378
rect 17390 4326 17392 4378
rect 17146 4324 17152 4326
rect 17208 4324 17232 4326
rect 17288 4324 17312 4326
rect 17368 4324 17392 4326
rect 17448 4324 17454 4326
rect 17146 4315 17454 4324
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 11900 3534 11928 4082
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8268 3292 8576 3301
rect 8268 3290 8274 3292
rect 8330 3290 8354 3292
rect 8410 3290 8434 3292
rect 8490 3290 8514 3292
rect 8570 3290 8576 3292
rect 8330 3238 8332 3290
rect 8512 3238 8514 3290
rect 8268 3236 8274 3238
rect 8330 3236 8354 3238
rect 8410 3236 8434 3238
rect 8490 3236 8514 3238
rect 8570 3236 8576 3238
rect 8268 3227 8576 3236
rect 12707 3292 13015 3301
rect 12707 3290 12713 3292
rect 12769 3290 12793 3292
rect 12849 3290 12873 3292
rect 12929 3290 12953 3292
rect 13009 3290 13015 3292
rect 12769 3238 12771 3290
rect 12951 3238 12953 3290
rect 12707 3236 12713 3238
rect 12769 3236 12793 3238
rect 12849 3236 12873 3238
rect 12929 3236 12953 3238
rect 13009 3236 13015 3238
rect 12707 3227 13015 3236
rect 17146 3292 17454 3301
rect 17146 3290 17152 3292
rect 17208 3290 17232 3292
rect 17288 3290 17312 3292
rect 17368 3290 17392 3292
rect 17448 3290 17454 3292
rect 17208 3238 17210 3290
rect 17390 3238 17392 3290
rect 17146 3236 17152 3238
rect 17208 3236 17232 3238
rect 17288 3236 17312 3238
rect 17368 3236 17392 3238
rect 17448 3236 17454 3238
rect 17146 3227 17454 3236
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5448 3052 5500 3058
rect 5368 3012 5448 3040
rect 5264 2994 5316 3000
rect 5448 2994 5500 3000
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 3829 2204 4137 2213
rect 3829 2202 3835 2204
rect 3891 2202 3915 2204
rect 3971 2202 3995 2204
rect 4051 2202 4075 2204
rect 4131 2202 4137 2204
rect 3891 2150 3893 2202
rect 4073 2150 4075 2202
rect 3829 2148 3835 2150
rect 3891 2148 3915 2150
rect 3971 2148 3995 2150
rect 4051 2148 4075 2150
rect 4131 2148 4137 2150
rect 3829 2139 4137 2148
rect 8268 2204 8576 2213
rect 8268 2202 8274 2204
rect 8330 2202 8354 2204
rect 8410 2202 8434 2204
rect 8490 2202 8514 2204
rect 8570 2202 8576 2204
rect 8330 2150 8332 2202
rect 8512 2150 8514 2202
rect 8268 2148 8274 2150
rect 8330 2148 8354 2150
rect 8410 2148 8434 2150
rect 8490 2148 8514 2150
rect 8570 2148 8576 2150
rect 8268 2139 8576 2148
rect 12707 2204 13015 2213
rect 12707 2202 12713 2204
rect 12769 2202 12793 2204
rect 12849 2202 12873 2204
rect 12929 2202 12953 2204
rect 13009 2202 13015 2204
rect 12769 2150 12771 2202
rect 12951 2150 12953 2202
rect 12707 2148 12713 2150
rect 12769 2148 12793 2150
rect 12849 2148 12873 2150
rect 12929 2148 12953 2150
rect 13009 2148 13015 2150
rect 12707 2139 13015 2148
rect 17146 2204 17454 2213
rect 17146 2202 17152 2204
rect 17208 2202 17232 2204
rect 17288 2202 17312 2204
rect 17368 2202 17392 2204
rect 17448 2202 17454 2204
rect 17208 2150 17210 2202
rect 17390 2150 17392 2202
rect 17146 2148 17152 2150
rect 17208 2148 17232 2150
rect 17288 2148 17312 2150
rect 17368 2148 17392 2150
rect 17448 2148 17454 2150
rect 17146 2139 17454 2148
<< via2 >>
rect 3835 7642 3891 7644
rect 3915 7642 3971 7644
rect 3995 7642 4051 7644
rect 4075 7642 4131 7644
rect 3835 7590 3881 7642
rect 3881 7590 3891 7642
rect 3915 7590 3945 7642
rect 3945 7590 3957 7642
rect 3957 7590 3971 7642
rect 3995 7590 4009 7642
rect 4009 7590 4021 7642
rect 4021 7590 4051 7642
rect 4075 7590 4085 7642
rect 4085 7590 4131 7642
rect 3835 7588 3891 7590
rect 3915 7588 3971 7590
rect 3995 7588 4051 7590
rect 4075 7588 4131 7590
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3835 6554 3891 6556
rect 3915 6554 3971 6556
rect 3995 6554 4051 6556
rect 4075 6554 4131 6556
rect 3835 6502 3881 6554
rect 3881 6502 3891 6554
rect 3915 6502 3945 6554
rect 3945 6502 3957 6554
rect 3957 6502 3971 6554
rect 3995 6502 4009 6554
rect 4009 6502 4021 6554
rect 4021 6502 4051 6554
rect 4075 6502 4085 6554
rect 4085 6502 4131 6554
rect 3835 6500 3891 6502
rect 3915 6500 3971 6502
rect 3995 6500 4051 6502
rect 4075 6500 4131 6502
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 3835 5466 3891 5468
rect 3915 5466 3971 5468
rect 3995 5466 4051 5468
rect 4075 5466 4131 5468
rect 3835 5414 3881 5466
rect 3881 5414 3891 5466
rect 3915 5414 3945 5466
rect 3945 5414 3957 5466
rect 3957 5414 3971 5466
rect 3995 5414 4009 5466
rect 4009 5414 4021 5466
rect 4021 5414 4051 5466
rect 4075 5414 4085 5466
rect 4085 5414 4131 5466
rect 3835 5412 3891 5414
rect 3915 5412 3971 5414
rect 3995 5412 4051 5414
rect 4075 5412 4131 5414
rect 4342 6860 4398 6896
rect 4342 6840 4344 6860
rect 4344 6840 4396 6860
rect 4396 6840 4398 6860
rect 4250 6568 4306 6624
rect 4342 5772 4398 5808
rect 4342 5752 4344 5772
rect 4344 5752 4396 5772
rect 4396 5752 4398 5772
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 3835 4378 3891 4380
rect 3915 4378 3971 4380
rect 3995 4378 4051 4380
rect 4075 4378 4131 4380
rect 3835 4326 3881 4378
rect 3881 4326 3891 4378
rect 3915 4326 3945 4378
rect 3945 4326 3957 4378
rect 3957 4326 3971 4378
rect 3995 4326 4009 4378
rect 4009 4326 4021 4378
rect 4021 4326 4051 4378
rect 4075 4326 4085 4378
rect 4085 4326 4131 4378
rect 3835 4324 3891 4326
rect 3915 4324 3971 4326
rect 3995 4324 4051 4326
rect 4075 4324 4131 4326
rect 5906 6840 5962 6896
rect 5722 6568 5778 6624
rect 5262 5752 5318 5808
rect 3835 3290 3891 3292
rect 3915 3290 3971 3292
rect 3995 3290 4051 3292
rect 4075 3290 4131 3292
rect 3835 3238 3881 3290
rect 3881 3238 3891 3290
rect 3915 3238 3945 3290
rect 3945 3238 3957 3290
rect 3957 3238 3971 3290
rect 3995 3238 4009 3290
rect 4009 3238 4021 3290
rect 4021 3238 4051 3290
rect 4075 3238 4085 3290
rect 4085 3238 4131 3290
rect 3835 3236 3891 3238
rect 3915 3236 3971 3238
rect 3995 3236 4051 3238
rect 4075 3236 4131 3238
rect 7286 5788 7288 5808
rect 7288 5788 7340 5808
rect 7340 5788 7342 5808
rect 7286 5752 7342 5788
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 8274 7642 8330 7644
rect 8354 7642 8410 7644
rect 8434 7642 8490 7644
rect 8514 7642 8570 7644
rect 8274 7590 8320 7642
rect 8320 7590 8330 7642
rect 8354 7590 8384 7642
rect 8384 7590 8396 7642
rect 8396 7590 8410 7642
rect 8434 7590 8448 7642
rect 8448 7590 8460 7642
rect 8460 7590 8490 7642
rect 8514 7590 8524 7642
rect 8524 7590 8570 7642
rect 8274 7588 8330 7590
rect 8354 7588 8410 7590
rect 8434 7588 8490 7590
rect 8514 7588 8570 7590
rect 8274 6554 8330 6556
rect 8354 6554 8410 6556
rect 8434 6554 8490 6556
rect 8514 6554 8570 6556
rect 8274 6502 8320 6554
rect 8320 6502 8330 6554
rect 8354 6502 8384 6554
rect 8384 6502 8396 6554
rect 8396 6502 8410 6554
rect 8434 6502 8448 6554
rect 8448 6502 8460 6554
rect 8460 6502 8490 6554
rect 8514 6502 8524 6554
rect 8524 6502 8570 6554
rect 8274 6500 8330 6502
rect 8354 6500 8410 6502
rect 8434 6500 8490 6502
rect 8514 6500 8570 6502
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 8274 5466 8330 5468
rect 8354 5466 8410 5468
rect 8434 5466 8490 5468
rect 8514 5466 8570 5468
rect 8274 5414 8320 5466
rect 8320 5414 8330 5466
rect 8354 5414 8384 5466
rect 8384 5414 8396 5466
rect 8396 5414 8410 5466
rect 8434 5414 8448 5466
rect 8448 5414 8460 5466
rect 8460 5414 8490 5466
rect 8514 5414 8524 5466
rect 8524 5414 8570 5466
rect 8274 5412 8330 5414
rect 8354 5412 8410 5414
rect 8434 5412 8490 5414
rect 8514 5412 8570 5414
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 8274 4378 8330 4380
rect 8354 4378 8410 4380
rect 8434 4378 8490 4380
rect 8514 4378 8570 4380
rect 8274 4326 8320 4378
rect 8320 4326 8330 4378
rect 8354 4326 8384 4378
rect 8384 4326 8396 4378
rect 8396 4326 8410 4378
rect 8434 4326 8448 4378
rect 8448 4326 8460 4378
rect 8460 4326 8490 4378
rect 8514 4326 8524 4378
rect 8524 4326 8570 4378
rect 8274 4324 8330 4326
rect 8354 4324 8410 4326
rect 8434 4324 8490 4326
rect 8514 4324 8570 4326
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 12713 7642 12769 7644
rect 12793 7642 12849 7644
rect 12873 7642 12929 7644
rect 12953 7642 13009 7644
rect 12713 7590 12759 7642
rect 12759 7590 12769 7642
rect 12793 7590 12823 7642
rect 12823 7590 12835 7642
rect 12835 7590 12849 7642
rect 12873 7590 12887 7642
rect 12887 7590 12899 7642
rect 12899 7590 12929 7642
rect 12953 7590 12963 7642
rect 12963 7590 13009 7642
rect 12713 7588 12769 7590
rect 12793 7588 12849 7590
rect 12873 7588 12929 7590
rect 12953 7588 13009 7590
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 12713 6554 12769 6556
rect 12793 6554 12849 6556
rect 12873 6554 12929 6556
rect 12953 6554 13009 6556
rect 12713 6502 12759 6554
rect 12759 6502 12769 6554
rect 12793 6502 12823 6554
rect 12823 6502 12835 6554
rect 12835 6502 12849 6554
rect 12873 6502 12887 6554
rect 12887 6502 12899 6554
rect 12899 6502 12929 6554
rect 12953 6502 12963 6554
rect 12963 6502 13009 6554
rect 12713 6500 12769 6502
rect 12793 6500 12849 6502
rect 12873 6500 12929 6502
rect 12953 6500 13009 6502
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 12713 5466 12769 5468
rect 12793 5466 12849 5468
rect 12873 5466 12929 5468
rect 12953 5466 13009 5468
rect 12713 5414 12759 5466
rect 12759 5414 12769 5466
rect 12793 5414 12823 5466
rect 12823 5414 12835 5466
rect 12835 5414 12849 5466
rect 12873 5414 12887 5466
rect 12887 5414 12899 5466
rect 12899 5414 12929 5466
rect 12953 5414 12963 5466
rect 12963 5414 13009 5466
rect 12713 5412 12769 5414
rect 12793 5412 12849 5414
rect 12873 5412 12929 5414
rect 12953 5412 13009 5414
rect 13726 6840 13782 6896
rect 17152 7642 17208 7644
rect 17232 7642 17288 7644
rect 17312 7642 17368 7644
rect 17392 7642 17448 7644
rect 17152 7590 17198 7642
rect 17198 7590 17208 7642
rect 17232 7590 17262 7642
rect 17262 7590 17274 7642
rect 17274 7590 17288 7642
rect 17312 7590 17326 7642
rect 17326 7590 17338 7642
rect 17338 7590 17368 7642
rect 17392 7590 17402 7642
rect 17402 7590 17448 7642
rect 17152 7588 17208 7590
rect 17232 7588 17288 7590
rect 17312 7588 17368 7590
rect 17392 7588 17448 7590
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 16854 6840 16910 6896
rect 17152 6554 17208 6556
rect 17232 6554 17288 6556
rect 17312 6554 17368 6556
rect 17392 6554 17448 6556
rect 17152 6502 17198 6554
rect 17198 6502 17208 6554
rect 17232 6502 17262 6554
rect 17262 6502 17274 6554
rect 17274 6502 17288 6554
rect 17312 6502 17326 6554
rect 17326 6502 17338 6554
rect 17338 6502 17368 6554
rect 17392 6502 17402 6554
rect 17402 6502 17448 6554
rect 17152 6500 17208 6502
rect 17232 6500 17288 6502
rect 17312 6500 17368 6502
rect 17392 6500 17448 6502
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 17152 5466 17208 5468
rect 17232 5466 17288 5468
rect 17312 5466 17368 5468
rect 17392 5466 17448 5468
rect 17152 5414 17198 5466
rect 17198 5414 17208 5466
rect 17232 5414 17262 5466
rect 17262 5414 17274 5466
rect 17274 5414 17288 5466
rect 17312 5414 17326 5466
rect 17326 5414 17338 5466
rect 17338 5414 17368 5466
rect 17392 5414 17402 5466
rect 17402 5414 17448 5466
rect 17152 5412 17208 5414
rect 17232 5412 17288 5414
rect 17312 5412 17368 5414
rect 17392 5412 17448 5414
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 12713 4378 12769 4380
rect 12793 4378 12849 4380
rect 12873 4378 12929 4380
rect 12953 4378 13009 4380
rect 12713 4326 12759 4378
rect 12759 4326 12769 4378
rect 12793 4326 12823 4378
rect 12823 4326 12835 4378
rect 12835 4326 12849 4378
rect 12873 4326 12887 4378
rect 12887 4326 12899 4378
rect 12899 4326 12929 4378
rect 12953 4326 12963 4378
rect 12963 4326 13009 4378
rect 12713 4324 12769 4326
rect 12793 4324 12849 4326
rect 12873 4324 12929 4326
rect 12953 4324 13009 4326
rect 17152 4378 17208 4380
rect 17232 4378 17288 4380
rect 17312 4378 17368 4380
rect 17392 4378 17448 4380
rect 17152 4326 17198 4378
rect 17198 4326 17208 4378
rect 17232 4326 17262 4378
rect 17262 4326 17274 4378
rect 17274 4326 17288 4378
rect 17312 4326 17326 4378
rect 17326 4326 17338 4378
rect 17338 4326 17368 4378
rect 17392 4326 17402 4378
rect 17402 4326 17448 4378
rect 17152 4324 17208 4326
rect 17232 4324 17288 4326
rect 17312 4324 17368 4326
rect 17392 4324 17448 4326
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 8274 3290 8330 3292
rect 8354 3290 8410 3292
rect 8434 3290 8490 3292
rect 8514 3290 8570 3292
rect 8274 3238 8320 3290
rect 8320 3238 8330 3290
rect 8354 3238 8384 3290
rect 8384 3238 8396 3290
rect 8396 3238 8410 3290
rect 8434 3238 8448 3290
rect 8448 3238 8460 3290
rect 8460 3238 8490 3290
rect 8514 3238 8524 3290
rect 8524 3238 8570 3290
rect 8274 3236 8330 3238
rect 8354 3236 8410 3238
rect 8434 3236 8490 3238
rect 8514 3236 8570 3238
rect 12713 3290 12769 3292
rect 12793 3290 12849 3292
rect 12873 3290 12929 3292
rect 12953 3290 13009 3292
rect 12713 3238 12759 3290
rect 12759 3238 12769 3290
rect 12793 3238 12823 3290
rect 12823 3238 12835 3290
rect 12835 3238 12849 3290
rect 12873 3238 12887 3290
rect 12887 3238 12899 3290
rect 12899 3238 12929 3290
rect 12953 3238 12963 3290
rect 12963 3238 13009 3290
rect 12713 3236 12769 3238
rect 12793 3236 12849 3238
rect 12873 3236 12929 3238
rect 12953 3236 13009 3238
rect 17152 3290 17208 3292
rect 17232 3290 17288 3292
rect 17312 3290 17368 3292
rect 17392 3290 17448 3292
rect 17152 3238 17198 3290
rect 17198 3238 17208 3290
rect 17232 3238 17262 3290
rect 17262 3238 17274 3290
rect 17274 3238 17288 3290
rect 17312 3238 17326 3290
rect 17326 3238 17338 3290
rect 17338 3238 17368 3290
rect 17392 3238 17402 3290
rect 17402 3238 17448 3290
rect 17152 3236 17208 3238
rect 17232 3236 17288 3238
rect 17312 3236 17368 3238
rect 17392 3236 17448 3238
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 3835 2202 3891 2204
rect 3915 2202 3971 2204
rect 3995 2202 4051 2204
rect 4075 2202 4131 2204
rect 3835 2150 3881 2202
rect 3881 2150 3891 2202
rect 3915 2150 3945 2202
rect 3945 2150 3957 2202
rect 3957 2150 3971 2202
rect 3995 2150 4009 2202
rect 4009 2150 4021 2202
rect 4021 2150 4051 2202
rect 4075 2150 4085 2202
rect 4085 2150 4131 2202
rect 3835 2148 3891 2150
rect 3915 2148 3971 2150
rect 3995 2148 4051 2150
rect 4075 2148 4131 2150
rect 8274 2202 8330 2204
rect 8354 2202 8410 2204
rect 8434 2202 8490 2204
rect 8514 2202 8570 2204
rect 8274 2150 8320 2202
rect 8320 2150 8330 2202
rect 8354 2150 8384 2202
rect 8384 2150 8396 2202
rect 8396 2150 8410 2202
rect 8434 2150 8448 2202
rect 8448 2150 8460 2202
rect 8460 2150 8490 2202
rect 8514 2150 8524 2202
rect 8524 2150 8570 2202
rect 8274 2148 8330 2150
rect 8354 2148 8410 2150
rect 8434 2148 8490 2150
rect 8514 2148 8570 2150
rect 12713 2202 12769 2204
rect 12793 2202 12849 2204
rect 12873 2202 12929 2204
rect 12953 2202 13009 2204
rect 12713 2150 12759 2202
rect 12759 2150 12769 2202
rect 12793 2150 12823 2202
rect 12823 2150 12835 2202
rect 12835 2150 12849 2202
rect 12873 2150 12887 2202
rect 12887 2150 12899 2202
rect 12899 2150 12929 2202
rect 12953 2150 12963 2202
rect 12963 2150 13009 2202
rect 12713 2148 12769 2150
rect 12793 2148 12849 2150
rect 12873 2148 12929 2150
rect 12953 2148 13009 2150
rect 17152 2202 17208 2204
rect 17232 2202 17288 2204
rect 17312 2202 17368 2204
rect 17392 2202 17448 2204
rect 17152 2150 17198 2202
rect 17198 2150 17208 2202
rect 17232 2150 17262 2202
rect 17262 2150 17274 2202
rect 17274 2150 17288 2202
rect 17312 2150 17326 2202
rect 17326 2150 17338 2202
rect 17338 2150 17368 2202
rect 17392 2150 17402 2202
rect 17402 2150 17448 2202
rect 17152 2148 17208 2150
rect 17232 2148 17288 2150
rect 17312 2148 17368 2150
rect 17392 2148 17448 2150
<< metal3 >>
rect 3825 7648 4141 7649
rect 3825 7584 3831 7648
rect 3895 7584 3911 7648
rect 3975 7584 3991 7648
rect 4055 7584 4071 7648
rect 4135 7584 4141 7648
rect 3825 7583 4141 7584
rect 8264 7648 8580 7649
rect 8264 7584 8270 7648
rect 8334 7584 8350 7648
rect 8414 7584 8430 7648
rect 8494 7584 8510 7648
rect 8574 7584 8580 7648
rect 8264 7583 8580 7584
rect 12703 7648 13019 7649
rect 12703 7584 12709 7648
rect 12773 7584 12789 7648
rect 12853 7584 12869 7648
rect 12933 7584 12949 7648
rect 13013 7584 13019 7648
rect 12703 7583 13019 7584
rect 17142 7648 17458 7649
rect 17142 7584 17148 7648
rect 17212 7584 17228 7648
rect 17292 7584 17308 7648
rect 17372 7584 17388 7648
rect 17452 7584 17458 7648
rect 17142 7583 17458 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 4337 6898 4403 6901
rect 5901 6898 5967 6901
rect 4337 6896 5967 6898
rect 4337 6840 4342 6896
rect 4398 6840 5906 6896
rect 5962 6840 5967 6896
rect 4337 6838 5967 6840
rect 4337 6835 4403 6838
rect 5901 6835 5967 6838
rect 13721 6898 13787 6901
rect 16849 6898 16915 6901
rect 13721 6896 16915 6898
rect 13721 6840 13726 6896
rect 13782 6840 16854 6896
rect 16910 6840 16915 6896
rect 13721 6838 16915 6840
rect 13721 6835 13787 6838
rect 16849 6835 16915 6838
rect 4245 6626 4311 6629
rect 5717 6626 5783 6629
rect 4245 6624 5783 6626
rect 4245 6568 4250 6624
rect 4306 6568 5722 6624
rect 5778 6568 5783 6624
rect 4245 6566 5783 6568
rect 4245 6563 4311 6566
rect 5717 6563 5783 6566
rect 3825 6560 4141 6561
rect 3825 6496 3831 6560
rect 3895 6496 3911 6560
rect 3975 6496 3991 6560
rect 4055 6496 4071 6560
rect 4135 6496 4141 6560
rect 3825 6495 4141 6496
rect 8264 6560 8580 6561
rect 8264 6496 8270 6560
rect 8334 6496 8350 6560
rect 8414 6496 8430 6560
rect 8494 6496 8510 6560
rect 8574 6496 8580 6560
rect 8264 6495 8580 6496
rect 12703 6560 13019 6561
rect 12703 6496 12709 6560
rect 12773 6496 12789 6560
rect 12853 6496 12869 6560
rect 12933 6496 12949 6560
rect 13013 6496 13019 6560
rect 12703 6495 13019 6496
rect 17142 6560 17458 6561
rect 17142 6496 17148 6560
rect 17212 6496 17228 6560
rect 17292 6496 17308 6560
rect 17372 6496 17388 6560
rect 17452 6496 17458 6560
rect 17142 6495 17458 6496
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 4337 5810 4403 5813
rect 5257 5810 5323 5813
rect 7281 5810 7347 5813
rect 4337 5808 7347 5810
rect 4337 5752 4342 5808
rect 4398 5752 5262 5808
rect 5318 5752 7286 5808
rect 7342 5752 7347 5808
rect 4337 5750 7347 5752
rect 4337 5747 4403 5750
rect 5257 5747 5323 5750
rect 7281 5747 7347 5750
rect 3825 5472 4141 5473
rect 3825 5408 3831 5472
rect 3895 5408 3911 5472
rect 3975 5408 3991 5472
rect 4055 5408 4071 5472
rect 4135 5408 4141 5472
rect 3825 5407 4141 5408
rect 8264 5472 8580 5473
rect 8264 5408 8270 5472
rect 8334 5408 8350 5472
rect 8414 5408 8430 5472
rect 8494 5408 8510 5472
rect 8574 5408 8580 5472
rect 8264 5407 8580 5408
rect 12703 5472 13019 5473
rect 12703 5408 12709 5472
rect 12773 5408 12789 5472
rect 12853 5408 12869 5472
rect 12933 5408 12949 5472
rect 13013 5408 13019 5472
rect 12703 5407 13019 5408
rect 17142 5472 17458 5473
rect 17142 5408 17148 5472
rect 17212 5408 17228 5472
rect 17292 5408 17308 5472
rect 17372 5408 17388 5472
rect 17452 5408 17458 5472
rect 17142 5407 17458 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 3825 4384 4141 4385
rect 3825 4320 3831 4384
rect 3895 4320 3911 4384
rect 3975 4320 3991 4384
rect 4055 4320 4071 4384
rect 4135 4320 4141 4384
rect 3825 4319 4141 4320
rect 8264 4384 8580 4385
rect 8264 4320 8270 4384
rect 8334 4320 8350 4384
rect 8414 4320 8430 4384
rect 8494 4320 8510 4384
rect 8574 4320 8580 4384
rect 8264 4319 8580 4320
rect 12703 4384 13019 4385
rect 12703 4320 12709 4384
rect 12773 4320 12789 4384
rect 12853 4320 12869 4384
rect 12933 4320 12949 4384
rect 13013 4320 13019 4384
rect 12703 4319 13019 4320
rect 17142 4384 17458 4385
rect 17142 4320 17148 4384
rect 17212 4320 17228 4384
rect 17292 4320 17308 4384
rect 17372 4320 17388 4384
rect 17452 4320 17458 4384
rect 17142 4319 17458 4320
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 3825 3296 4141 3297
rect 3825 3232 3831 3296
rect 3895 3232 3911 3296
rect 3975 3232 3991 3296
rect 4055 3232 4071 3296
rect 4135 3232 4141 3296
rect 3825 3231 4141 3232
rect 8264 3296 8580 3297
rect 8264 3232 8270 3296
rect 8334 3232 8350 3296
rect 8414 3232 8430 3296
rect 8494 3232 8510 3296
rect 8574 3232 8580 3296
rect 8264 3231 8580 3232
rect 12703 3296 13019 3297
rect 12703 3232 12709 3296
rect 12773 3232 12789 3296
rect 12853 3232 12869 3296
rect 12933 3232 12949 3296
rect 13013 3232 13019 3296
rect 12703 3231 13019 3232
rect 17142 3296 17458 3297
rect 17142 3232 17148 3296
rect 17212 3232 17228 3296
rect 17292 3232 17308 3296
rect 17372 3232 17388 3296
rect 17452 3232 17458 3296
rect 17142 3231 17458 3232
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 3825 2208 4141 2209
rect 3825 2144 3831 2208
rect 3895 2144 3911 2208
rect 3975 2144 3991 2208
rect 4055 2144 4071 2208
rect 4135 2144 4141 2208
rect 3825 2143 4141 2144
rect 8264 2208 8580 2209
rect 8264 2144 8270 2208
rect 8334 2144 8350 2208
rect 8414 2144 8430 2208
rect 8494 2144 8510 2208
rect 8574 2144 8580 2208
rect 8264 2143 8580 2144
rect 12703 2208 13019 2209
rect 12703 2144 12709 2208
rect 12773 2144 12789 2208
rect 12853 2144 12869 2208
rect 12933 2144 12949 2208
rect 13013 2144 13019 2208
rect 12703 2143 13019 2144
rect 17142 2208 17458 2209
rect 17142 2144 17148 2208
rect 17212 2144 17228 2208
rect 17292 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17458 2208
rect 17142 2143 17458 2144
<< via3 >>
rect 3831 7644 3895 7648
rect 3831 7588 3835 7644
rect 3835 7588 3891 7644
rect 3891 7588 3895 7644
rect 3831 7584 3895 7588
rect 3911 7644 3975 7648
rect 3911 7588 3915 7644
rect 3915 7588 3971 7644
rect 3971 7588 3975 7644
rect 3911 7584 3975 7588
rect 3991 7644 4055 7648
rect 3991 7588 3995 7644
rect 3995 7588 4051 7644
rect 4051 7588 4055 7644
rect 3991 7584 4055 7588
rect 4071 7644 4135 7648
rect 4071 7588 4075 7644
rect 4075 7588 4131 7644
rect 4131 7588 4135 7644
rect 4071 7584 4135 7588
rect 8270 7644 8334 7648
rect 8270 7588 8274 7644
rect 8274 7588 8330 7644
rect 8330 7588 8334 7644
rect 8270 7584 8334 7588
rect 8350 7644 8414 7648
rect 8350 7588 8354 7644
rect 8354 7588 8410 7644
rect 8410 7588 8414 7644
rect 8350 7584 8414 7588
rect 8430 7644 8494 7648
rect 8430 7588 8434 7644
rect 8434 7588 8490 7644
rect 8490 7588 8494 7644
rect 8430 7584 8494 7588
rect 8510 7644 8574 7648
rect 8510 7588 8514 7644
rect 8514 7588 8570 7644
rect 8570 7588 8574 7644
rect 8510 7584 8574 7588
rect 12709 7644 12773 7648
rect 12709 7588 12713 7644
rect 12713 7588 12769 7644
rect 12769 7588 12773 7644
rect 12709 7584 12773 7588
rect 12789 7644 12853 7648
rect 12789 7588 12793 7644
rect 12793 7588 12849 7644
rect 12849 7588 12853 7644
rect 12789 7584 12853 7588
rect 12869 7644 12933 7648
rect 12869 7588 12873 7644
rect 12873 7588 12929 7644
rect 12929 7588 12933 7644
rect 12869 7584 12933 7588
rect 12949 7644 13013 7648
rect 12949 7588 12953 7644
rect 12953 7588 13009 7644
rect 13009 7588 13013 7644
rect 12949 7584 13013 7588
rect 17148 7644 17212 7648
rect 17148 7588 17152 7644
rect 17152 7588 17208 7644
rect 17208 7588 17212 7644
rect 17148 7584 17212 7588
rect 17228 7644 17292 7648
rect 17228 7588 17232 7644
rect 17232 7588 17288 7644
rect 17288 7588 17292 7644
rect 17228 7584 17292 7588
rect 17308 7644 17372 7648
rect 17308 7588 17312 7644
rect 17312 7588 17368 7644
rect 17368 7588 17372 7644
rect 17308 7584 17372 7588
rect 17388 7644 17452 7648
rect 17388 7588 17392 7644
rect 17392 7588 17448 7644
rect 17448 7588 17452 7644
rect 17388 7584 17452 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 3831 6556 3895 6560
rect 3831 6500 3835 6556
rect 3835 6500 3891 6556
rect 3891 6500 3895 6556
rect 3831 6496 3895 6500
rect 3911 6556 3975 6560
rect 3911 6500 3915 6556
rect 3915 6500 3971 6556
rect 3971 6500 3975 6556
rect 3911 6496 3975 6500
rect 3991 6556 4055 6560
rect 3991 6500 3995 6556
rect 3995 6500 4051 6556
rect 4051 6500 4055 6556
rect 3991 6496 4055 6500
rect 4071 6556 4135 6560
rect 4071 6500 4075 6556
rect 4075 6500 4131 6556
rect 4131 6500 4135 6556
rect 4071 6496 4135 6500
rect 8270 6556 8334 6560
rect 8270 6500 8274 6556
rect 8274 6500 8330 6556
rect 8330 6500 8334 6556
rect 8270 6496 8334 6500
rect 8350 6556 8414 6560
rect 8350 6500 8354 6556
rect 8354 6500 8410 6556
rect 8410 6500 8414 6556
rect 8350 6496 8414 6500
rect 8430 6556 8494 6560
rect 8430 6500 8434 6556
rect 8434 6500 8490 6556
rect 8490 6500 8494 6556
rect 8430 6496 8494 6500
rect 8510 6556 8574 6560
rect 8510 6500 8514 6556
rect 8514 6500 8570 6556
rect 8570 6500 8574 6556
rect 8510 6496 8574 6500
rect 12709 6556 12773 6560
rect 12709 6500 12713 6556
rect 12713 6500 12769 6556
rect 12769 6500 12773 6556
rect 12709 6496 12773 6500
rect 12789 6556 12853 6560
rect 12789 6500 12793 6556
rect 12793 6500 12849 6556
rect 12849 6500 12853 6556
rect 12789 6496 12853 6500
rect 12869 6556 12933 6560
rect 12869 6500 12873 6556
rect 12873 6500 12929 6556
rect 12929 6500 12933 6556
rect 12869 6496 12933 6500
rect 12949 6556 13013 6560
rect 12949 6500 12953 6556
rect 12953 6500 13009 6556
rect 13009 6500 13013 6556
rect 12949 6496 13013 6500
rect 17148 6556 17212 6560
rect 17148 6500 17152 6556
rect 17152 6500 17208 6556
rect 17208 6500 17212 6556
rect 17148 6496 17212 6500
rect 17228 6556 17292 6560
rect 17228 6500 17232 6556
rect 17232 6500 17288 6556
rect 17288 6500 17292 6556
rect 17228 6496 17292 6500
rect 17308 6556 17372 6560
rect 17308 6500 17312 6556
rect 17312 6500 17368 6556
rect 17368 6500 17372 6556
rect 17308 6496 17372 6500
rect 17388 6556 17452 6560
rect 17388 6500 17392 6556
rect 17392 6500 17448 6556
rect 17448 6500 17452 6556
rect 17388 6496 17452 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 3831 5468 3895 5472
rect 3831 5412 3835 5468
rect 3835 5412 3891 5468
rect 3891 5412 3895 5468
rect 3831 5408 3895 5412
rect 3911 5468 3975 5472
rect 3911 5412 3915 5468
rect 3915 5412 3971 5468
rect 3971 5412 3975 5468
rect 3911 5408 3975 5412
rect 3991 5468 4055 5472
rect 3991 5412 3995 5468
rect 3995 5412 4051 5468
rect 4051 5412 4055 5468
rect 3991 5408 4055 5412
rect 4071 5468 4135 5472
rect 4071 5412 4075 5468
rect 4075 5412 4131 5468
rect 4131 5412 4135 5468
rect 4071 5408 4135 5412
rect 8270 5468 8334 5472
rect 8270 5412 8274 5468
rect 8274 5412 8330 5468
rect 8330 5412 8334 5468
rect 8270 5408 8334 5412
rect 8350 5468 8414 5472
rect 8350 5412 8354 5468
rect 8354 5412 8410 5468
rect 8410 5412 8414 5468
rect 8350 5408 8414 5412
rect 8430 5468 8494 5472
rect 8430 5412 8434 5468
rect 8434 5412 8490 5468
rect 8490 5412 8494 5468
rect 8430 5408 8494 5412
rect 8510 5468 8574 5472
rect 8510 5412 8514 5468
rect 8514 5412 8570 5468
rect 8570 5412 8574 5468
rect 8510 5408 8574 5412
rect 12709 5468 12773 5472
rect 12709 5412 12713 5468
rect 12713 5412 12769 5468
rect 12769 5412 12773 5468
rect 12709 5408 12773 5412
rect 12789 5468 12853 5472
rect 12789 5412 12793 5468
rect 12793 5412 12849 5468
rect 12849 5412 12853 5468
rect 12789 5408 12853 5412
rect 12869 5468 12933 5472
rect 12869 5412 12873 5468
rect 12873 5412 12929 5468
rect 12929 5412 12933 5468
rect 12869 5408 12933 5412
rect 12949 5468 13013 5472
rect 12949 5412 12953 5468
rect 12953 5412 13009 5468
rect 13009 5412 13013 5468
rect 12949 5408 13013 5412
rect 17148 5468 17212 5472
rect 17148 5412 17152 5468
rect 17152 5412 17208 5468
rect 17208 5412 17212 5468
rect 17148 5408 17212 5412
rect 17228 5468 17292 5472
rect 17228 5412 17232 5468
rect 17232 5412 17288 5468
rect 17288 5412 17292 5468
rect 17228 5408 17292 5412
rect 17308 5468 17372 5472
rect 17308 5412 17312 5468
rect 17312 5412 17368 5468
rect 17368 5412 17372 5468
rect 17308 5408 17372 5412
rect 17388 5468 17452 5472
rect 17388 5412 17392 5468
rect 17392 5412 17448 5468
rect 17448 5412 17452 5468
rect 17388 5408 17452 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 3831 4380 3895 4384
rect 3831 4324 3835 4380
rect 3835 4324 3891 4380
rect 3891 4324 3895 4380
rect 3831 4320 3895 4324
rect 3911 4380 3975 4384
rect 3911 4324 3915 4380
rect 3915 4324 3971 4380
rect 3971 4324 3975 4380
rect 3911 4320 3975 4324
rect 3991 4380 4055 4384
rect 3991 4324 3995 4380
rect 3995 4324 4051 4380
rect 4051 4324 4055 4380
rect 3991 4320 4055 4324
rect 4071 4380 4135 4384
rect 4071 4324 4075 4380
rect 4075 4324 4131 4380
rect 4131 4324 4135 4380
rect 4071 4320 4135 4324
rect 8270 4380 8334 4384
rect 8270 4324 8274 4380
rect 8274 4324 8330 4380
rect 8330 4324 8334 4380
rect 8270 4320 8334 4324
rect 8350 4380 8414 4384
rect 8350 4324 8354 4380
rect 8354 4324 8410 4380
rect 8410 4324 8414 4380
rect 8350 4320 8414 4324
rect 8430 4380 8494 4384
rect 8430 4324 8434 4380
rect 8434 4324 8490 4380
rect 8490 4324 8494 4380
rect 8430 4320 8494 4324
rect 8510 4380 8574 4384
rect 8510 4324 8514 4380
rect 8514 4324 8570 4380
rect 8570 4324 8574 4380
rect 8510 4320 8574 4324
rect 12709 4380 12773 4384
rect 12709 4324 12713 4380
rect 12713 4324 12769 4380
rect 12769 4324 12773 4380
rect 12709 4320 12773 4324
rect 12789 4380 12853 4384
rect 12789 4324 12793 4380
rect 12793 4324 12849 4380
rect 12849 4324 12853 4380
rect 12789 4320 12853 4324
rect 12869 4380 12933 4384
rect 12869 4324 12873 4380
rect 12873 4324 12929 4380
rect 12929 4324 12933 4380
rect 12869 4320 12933 4324
rect 12949 4380 13013 4384
rect 12949 4324 12953 4380
rect 12953 4324 13009 4380
rect 13009 4324 13013 4380
rect 12949 4320 13013 4324
rect 17148 4380 17212 4384
rect 17148 4324 17152 4380
rect 17152 4324 17208 4380
rect 17208 4324 17212 4380
rect 17148 4320 17212 4324
rect 17228 4380 17292 4384
rect 17228 4324 17232 4380
rect 17232 4324 17288 4380
rect 17288 4324 17292 4380
rect 17228 4320 17292 4324
rect 17308 4380 17372 4384
rect 17308 4324 17312 4380
rect 17312 4324 17368 4380
rect 17368 4324 17372 4380
rect 17308 4320 17372 4324
rect 17388 4380 17452 4384
rect 17388 4324 17392 4380
rect 17392 4324 17448 4380
rect 17448 4324 17452 4380
rect 17388 4320 17452 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 3831 3292 3895 3296
rect 3831 3236 3835 3292
rect 3835 3236 3891 3292
rect 3891 3236 3895 3292
rect 3831 3232 3895 3236
rect 3911 3292 3975 3296
rect 3911 3236 3915 3292
rect 3915 3236 3971 3292
rect 3971 3236 3975 3292
rect 3911 3232 3975 3236
rect 3991 3292 4055 3296
rect 3991 3236 3995 3292
rect 3995 3236 4051 3292
rect 4051 3236 4055 3292
rect 3991 3232 4055 3236
rect 4071 3292 4135 3296
rect 4071 3236 4075 3292
rect 4075 3236 4131 3292
rect 4131 3236 4135 3292
rect 4071 3232 4135 3236
rect 8270 3292 8334 3296
rect 8270 3236 8274 3292
rect 8274 3236 8330 3292
rect 8330 3236 8334 3292
rect 8270 3232 8334 3236
rect 8350 3292 8414 3296
rect 8350 3236 8354 3292
rect 8354 3236 8410 3292
rect 8410 3236 8414 3292
rect 8350 3232 8414 3236
rect 8430 3292 8494 3296
rect 8430 3236 8434 3292
rect 8434 3236 8490 3292
rect 8490 3236 8494 3292
rect 8430 3232 8494 3236
rect 8510 3292 8574 3296
rect 8510 3236 8514 3292
rect 8514 3236 8570 3292
rect 8570 3236 8574 3292
rect 8510 3232 8574 3236
rect 12709 3292 12773 3296
rect 12709 3236 12713 3292
rect 12713 3236 12769 3292
rect 12769 3236 12773 3292
rect 12709 3232 12773 3236
rect 12789 3292 12853 3296
rect 12789 3236 12793 3292
rect 12793 3236 12849 3292
rect 12849 3236 12853 3292
rect 12789 3232 12853 3236
rect 12869 3292 12933 3296
rect 12869 3236 12873 3292
rect 12873 3236 12929 3292
rect 12929 3236 12933 3292
rect 12869 3232 12933 3236
rect 12949 3292 13013 3296
rect 12949 3236 12953 3292
rect 12953 3236 13009 3292
rect 13009 3236 13013 3292
rect 12949 3232 13013 3236
rect 17148 3292 17212 3296
rect 17148 3236 17152 3292
rect 17152 3236 17208 3292
rect 17208 3236 17212 3292
rect 17148 3232 17212 3236
rect 17228 3292 17292 3296
rect 17228 3236 17232 3292
rect 17232 3236 17288 3292
rect 17288 3236 17292 3292
rect 17228 3232 17292 3236
rect 17308 3292 17372 3296
rect 17308 3236 17312 3292
rect 17312 3236 17368 3292
rect 17368 3236 17372 3292
rect 17308 3232 17372 3236
rect 17388 3292 17452 3296
rect 17388 3236 17392 3292
rect 17392 3236 17448 3292
rect 17448 3236 17452 3292
rect 17388 3232 17452 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 3831 2204 3895 2208
rect 3831 2148 3835 2204
rect 3835 2148 3891 2204
rect 3891 2148 3895 2204
rect 3831 2144 3895 2148
rect 3911 2204 3975 2208
rect 3911 2148 3915 2204
rect 3915 2148 3971 2204
rect 3971 2148 3975 2204
rect 3911 2144 3975 2148
rect 3991 2204 4055 2208
rect 3991 2148 3995 2204
rect 3995 2148 4051 2204
rect 4051 2148 4055 2204
rect 3991 2144 4055 2148
rect 4071 2204 4135 2208
rect 4071 2148 4075 2204
rect 4075 2148 4131 2204
rect 4131 2148 4135 2204
rect 4071 2144 4135 2148
rect 8270 2204 8334 2208
rect 8270 2148 8274 2204
rect 8274 2148 8330 2204
rect 8330 2148 8334 2204
rect 8270 2144 8334 2148
rect 8350 2204 8414 2208
rect 8350 2148 8354 2204
rect 8354 2148 8410 2204
rect 8410 2148 8414 2204
rect 8350 2144 8414 2148
rect 8430 2204 8494 2208
rect 8430 2148 8434 2204
rect 8434 2148 8490 2204
rect 8490 2148 8494 2204
rect 8430 2144 8494 2148
rect 8510 2204 8574 2208
rect 8510 2148 8514 2204
rect 8514 2148 8570 2204
rect 8570 2148 8574 2204
rect 8510 2144 8574 2148
rect 12709 2204 12773 2208
rect 12709 2148 12713 2204
rect 12713 2148 12769 2204
rect 12769 2148 12773 2204
rect 12709 2144 12773 2148
rect 12789 2204 12853 2208
rect 12789 2148 12793 2204
rect 12793 2148 12849 2204
rect 12849 2148 12853 2204
rect 12789 2144 12853 2148
rect 12869 2204 12933 2208
rect 12869 2148 12873 2204
rect 12873 2148 12929 2204
rect 12929 2148 12933 2204
rect 12869 2144 12933 2148
rect 12949 2204 13013 2208
rect 12949 2148 12953 2204
rect 12953 2148 13009 2204
rect 13009 2148 13013 2204
rect 12949 2144 13013 2148
rect 17148 2204 17212 2208
rect 17148 2148 17152 2204
rect 17152 2148 17208 2204
rect 17208 2148 17212 2204
rect 17148 2144 17212 2148
rect 17228 2204 17292 2208
rect 17228 2148 17232 2204
rect 17232 2148 17288 2204
rect 17288 2148 17292 2204
rect 17228 2144 17292 2148
rect 17308 2204 17372 2208
rect 17308 2148 17312 2204
rect 17312 2148 17368 2204
rect 17368 2148 17372 2204
rect 17308 2144 17372 2148
rect 17388 2204 17452 2208
rect 17388 2148 17392 2204
rect 17392 2148 17448 2204
rect 17448 2148 17452 2204
rect 17388 2144 17452 2148
<< metal4 >>
rect 3823 7710 4143 7752
rect 3163 7104 3483 7664
rect 3163 7040 3171 7104
rect 3235 7050 3251 7104
rect 3315 7050 3331 7104
rect 3395 7050 3411 7104
rect 3475 7040 3483 7104
rect 3163 6814 3205 7040
rect 3441 6814 3483 7040
rect 3163 6016 3483 6814
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 5691 3483 5952
rect 3163 5455 3205 5691
rect 3441 5455 3483 5691
rect 3163 4928 3483 5455
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 4332 3483 4864
rect 3163 4096 3205 4332
rect 3441 4096 3483 4332
rect 3163 3840 3483 4096
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2973 3483 3776
rect 3163 2752 3205 2973
rect 3441 2752 3483 2973
rect 3163 2688 3171 2752
rect 3235 2688 3251 2737
rect 3315 2688 3331 2737
rect 3395 2688 3411 2737
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 3823 7648 3865 7710
rect 4101 7648 4143 7710
rect 8262 7710 8582 7752
rect 3823 7584 3831 7648
rect 4135 7584 4143 7648
rect 3823 7474 3865 7584
rect 4101 7474 4143 7584
rect 3823 6560 4143 7474
rect 3823 6496 3831 6560
rect 3895 6496 3911 6560
rect 3975 6496 3991 6560
rect 4055 6496 4071 6560
rect 4135 6496 4143 6560
rect 3823 6351 4143 6496
rect 3823 6115 3865 6351
rect 4101 6115 4143 6351
rect 3823 5472 4143 6115
rect 3823 5408 3831 5472
rect 3895 5408 3911 5472
rect 3975 5408 3991 5472
rect 4055 5408 4071 5472
rect 4135 5408 4143 5472
rect 3823 4992 4143 5408
rect 3823 4756 3865 4992
rect 4101 4756 4143 4992
rect 3823 4384 4143 4756
rect 3823 4320 3831 4384
rect 3895 4320 3911 4384
rect 3975 4320 3991 4384
rect 4055 4320 4071 4384
rect 4135 4320 4143 4384
rect 3823 3633 4143 4320
rect 3823 3397 3865 3633
rect 4101 3397 4143 3633
rect 3823 3296 4143 3397
rect 3823 3232 3831 3296
rect 3895 3232 3911 3296
rect 3975 3232 3991 3296
rect 4055 3232 4071 3296
rect 4135 3232 4143 3296
rect 3823 2208 4143 3232
rect 3823 2144 3831 2208
rect 3895 2144 3911 2208
rect 3975 2144 3991 2208
rect 4055 2144 4071 2208
rect 4135 2144 4143 2208
rect 3823 2128 4143 2144
rect 7602 7104 7922 7664
rect 7602 7040 7610 7104
rect 7674 7050 7690 7104
rect 7754 7050 7770 7104
rect 7834 7050 7850 7104
rect 7914 7040 7922 7104
rect 7602 6814 7644 7040
rect 7880 6814 7922 7040
rect 7602 6016 7922 6814
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 5691 7922 5952
rect 7602 5455 7644 5691
rect 7880 5455 7922 5691
rect 7602 4928 7922 5455
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 4332 7922 4864
rect 7602 4096 7644 4332
rect 7880 4096 7922 4332
rect 7602 3840 7922 4096
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2973 7922 3776
rect 7602 2752 7644 2973
rect 7880 2752 7922 2973
rect 7602 2688 7610 2752
rect 7674 2688 7690 2737
rect 7754 2688 7770 2737
rect 7834 2688 7850 2737
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 8262 7648 8304 7710
rect 8540 7648 8582 7710
rect 12701 7710 13021 7752
rect 8262 7584 8270 7648
rect 8574 7584 8582 7648
rect 8262 7474 8304 7584
rect 8540 7474 8582 7584
rect 8262 6560 8582 7474
rect 8262 6496 8270 6560
rect 8334 6496 8350 6560
rect 8414 6496 8430 6560
rect 8494 6496 8510 6560
rect 8574 6496 8582 6560
rect 8262 6351 8582 6496
rect 8262 6115 8304 6351
rect 8540 6115 8582 6351
rect 8262 5472 8582 6115
rect 8262 5408 8270 5472
rect 8334 5408 8350 5472
rect 8414 5408 8430 5472
rect 8494 5408 8510 5472
rect 8574 5408 8582 5472
rect 8262 4992 8582 5408
rect 8262 4756 8304 4992
rect 8540 4756 8582 4992
rect 8262 4384 8582 4756
rect 8262 4320 8270 4384
rect 8334 4320 8350 4384
rect 8414 4320 8430 4384
rect 8494 4320 8510 4384
rect 8574 4320 8582 4384
rect 8262 3633 8582 4320
rect 8262 3397 8304 3633
rect 8540 3397 8582 3633
rect 8262 3296 8582 3397
rect 8262 3232 8270 3296
rect 8334 3232 8350 3296
rect 8414 3232 8430 3296
rect 8494 3232 8510 3296
rect 8574 3232 8582 3296
rect 8262 2208 8582 3232
rect 8262 2144 8270 2208
rect 8334 2144 8350 2208
rect 8414 2144 8430 2208
rect 8494 2144 8510 2208
rect 8574 2144 8582 2208
rect 8262 2128 8582 2144
rect 12041 7104 12361 7664
rect 12041 7040 12049 7104
rect 12113 7050 12129 7104
rect 12193 7050 12209 7104
rect 12273 7050 12289 7104
rect 12353 7040 12361 7104
rect 12041 6814 12083 7040
rect 12319 6814 12361 7040
rect 12041 6016 12361 6814
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 5691 12361 5952
rect 12041 5455 12083 5691
rect 12319 5455 12361 5691
rect 12041 4928 12361 5455
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 4332 12361 4864
rect 12041 4096 12083 4332
rect 12319 4096 12361 4332
rect 12041 3840 12361 4096
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2973 12361 3776
rect 12041 2752 12083 2973
rect 12319 2752 12361 2973
rect 12041 2688 12049 2752
rect 12113 2688 12129 2737
rect 12193 2688 12209 2737
rect 12273 2688 12289 2737
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 12701 7648 12743 7710
rect 12979 7648 13021 7710
rect 17140 7710 17460 7752
rect 12701 7584 12709 7648
rect 13013 7584 13021 7648
rect 12701 7474 12743 7584
rect 12979 7474 13021 7584
rect 12701 6560 13021 7474
rect 12701 6496 12709 6560
rect 12773 6496 12789 6560
rect 12853 6496 12869 6560
rect 12933 6496 12949 6560
rect 13013 6496 13021 6560
rect 12701 6351 13021 6496
rect 12701 6115 12743 6351
rect 12979 6115 13021 6351
rect 12701 5472 13021 6115
rect 12701 5408 12709 5472
rect 12773 5408 12789 5472
rect 12853 5408 12869 5472
rect 12933 5408 12949 5472
rect 13013 5408 13021 5472
rect 12701 4992 13021 5408
rect 12701 4756 12743 4992
rect 12979 4756 13021 4992
rect 12701 4384 13021 4756
rect 12701 4320 12709 4384
rect 12773 4320 12789 4384
rect 12853 4320 12869 4384
rect 12933 4320 12949 4384
rect 13013 4320 13021 4384
rect 12701 3633 13021 4320
rect 12701 3397 12743 3633
rect 12979 3397 13021 3633
rect 12701 3296 13021 3397
rect 12701 3232 12709 3296
rect 12773 3232 12789 3296
rect 12853 3232 12869 3296
rect 12933 3232 12949 3296
rect 13013 3232 13021 3296
rect 12701 2208 13021 3232
rect 12701 2144 12709 2208
rect 12773 2144 12789 2208
rect 12853 2144 12869 2208
rect 12933 2144 12949 2208
rect 13013 2144 13021 2208
rect 12701 2128 13021 2144
rect 16480 7104 16800 7664
rect 16480 7040 16488 7104
rect 16552 7050 16568 7104
rect 16632 7050 16648 7104
rect 16712 7050 16728 7104
rect 16792 7040 16800 7104
rect 16480 6814 16522 7040
rect 16758 6814 16800 7040
rect 16480 6016 16800 6814
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 5691 16800 5952
rect 16480 5455 16522 5691
rect 16758 5455 16800 5691
rect 16480 4928 16800 5455
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 4332 16800 4864
rect 16480 4096 16522 4332
rect 16758 4096 16800 4332
rect 16480 3840 16800 4096
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2973 16800 3776
rect 16480 2752 16522 2973
rect 16758 2752 16800 2973
rect 16480 2688 16488 2752
rect 16552 2688 16568 2737
rect 16632 2688 16648 2737
rect 16712 2688 16728 2737
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 17140 7648 17182 7710
rect 17418 7648 17460 7710
rect 17140 7584 17148 7648
rect 17452 7584 17460 7648
rect 17140 7474 17182 7584
rect 17418 7474 17460 7584
rect 17140 6560 17460 7474
rect 17140 6496 17148 6560
rect 17212 6496 17228 6560
rect 17292 6496 17308 6560
rect 17372 6496 17388 6560
rect 17452 6496 17460 6560
rect 17140 6351 17460 6496
rect 17140 6115 17182 6351
rect 17418 6115 17460 6351
rect 17140 5472 17460 6115
rect 17140 5408 17148 5472
rect 17212 5408 17228 5472
rect 17292 5408 17308 5472
rect 17372 5408 17388 5472
rect 17452 5408 17460 5472
rect 17140 4992 17460 5408
rect 17140 4756 17182 4992
rect 17418 4756 17460 4992
rect 17140 4384 17460 4756
rect 17140 4320 17148 4384
rect 17212 4320 17228 4384
rect 17292 4320 17308 4384
rect 17372 4320 17388 4384
rect 17452 4320 17460 4384
rect 17140 3633 17460 4320
rect 17140 3397 17182 3633
rect 17418 3397 17460 3633
rect 17140 3296 17460 3397
rect 17140 3232 17148 3296
rect 17212 3232 17228 3296
rect 17292 3232 17308 3296
rect 17372 3232 17388 3296
rect 17452 3232 17460 3296
rect 17140 2208 17460 3232
rect 17140 2144 17148 2208
rect 17212 2144 17228 2208
rect 17292 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17460 2208
rect 17140 2128 17460 2144
<< via4 >>
rect 3205 7040 3235 7050
rect 3235 7040 3251 7050
rect 3251 7040 3315 7050
rect 3315 7040 3331 7050
rect 3331 7040 3395 7050
rect 3395 7040 3411 7050
rect 3411 7040 3441 7050
rect 3205 6814 3441 7040
rect 3205 5455 3441 5691
rect 3205 4096 3441 4332
rect 3205 2752 3441 2973
rect 3205 2737 3235 2752
rect 3235 2737 3251 2752
rect 3251 2737 3315 2752
rect 3315 2737 3331 2752
rect 3331 2737 3395 2752
rect 3395 2737 3411 2752
rect 3411 2737 3441 2752
rect 3865 7648 4101 7710
rect 3865 7584 3895 7648
rect 3895 7584 3911 7648
rect 3911 7584 3975 7648
rect 3975 7584 3991 7648
rect 3991 7584 4055 7648
rect 4055 7584 4071 7648
rect 4071 7584 4101 7648
rect 3865 7474 4101 7584
rect 3865 6115 4101 6351
rect 3865 4756 4101 4992
rect 3865 3397 4101 3633
rect 7644 7040 7674 7050
rect 7674 7040 7690 7050
rect 7690 7040 7754 7050
rect 7754 7040 7770 7050
rect 7770 7040 7834 7050
rect 7834 7040 7850 7050
rect 7850 7040 7880 7050
rect 7644 6814 7880 7040
rect 7644 5455 7880 5691
rect 7644 4096 7880 4332
rect 7644 2752 7880 2973
rect 7644 2737 7674 2752
rect 7674 2737 7690 2752
rect 7690 2737 7754 2752
rect 7754 2737 7770 2752
rect 7770 2737 7834 2752
rect 7834 2737 7850 2752
rect 7850 2737 7880 2752
rect 8304 7648 8540 7710
rect 8304 7584 8334 7648
rect 8334 7584 8350 7648
rect 8350 7584 8414 7648
rect 8414 7584 8430 7648
rect 8430 7584 8494 7648
rect 8494 7584 8510 7648
rect 8510 7584 8540 7648
rect 8304 7474 8540 7584
rect 8304 6115 8540 6351
rect 8304 4756 8540 4992
rect 8304 3397 8540 3633
rect 12083 7040 12113 7050
rect 12113 7040 12129 7050
rect 12129 7040 12193 7050
rect 12193 7040 12209 7050
rect 12209 7040 12273 7050
rect 12273 7040 12289 7050
rect 12289 7040 12319 7050
rect 12083 6814 12319 7040
rect 12083 5455 12319 5691
rect 12083 4096 12319 4332
rect 12083 2752 12319 2973
rect 12083 2737 12113 2752
rect 12113 2737 12129 2752
rect 12129 2737 12193 2752
rect 12193 2737 12209 2752
rect 12209 2737 12273 2752
rect 12273 2737 12289 2752
rect 12289 2737 12319 2752
rect 12743 7648 12979 7710
rect 12743 7584 12773 7648
rect 12773 7584 12789 7648
rect 12789 7584 12853 7648
rect 12853 7584 12869 7648
rect 12869 7584 12933 7648
rect 12933 7584 12949 7648
rect 12949 7584 12979 7648
rect 12743 7474 12979 7584
rect 12743 6115 12979 6351
rect 12743 4756 12979 4992
rect 12743 3397 12979 3633
rect 16522 7040 16552 7050
rect 16552 7040 16568 7050
rect 16568 7040 16632 7050
rect 16632 7040 16648 7050
rect 16648 7040 16712 7050
rect 16712 7040 16728 7050
rect 16728 7040 16758 7050
rect 16522 6814 16758 7040
rect 16522 5455 16758 5691
rect 16522 4096 16758 4332
rect 16522 2752 16758 2973
rect 16522 2737 16552 2752
rect 16552 2737 16568 2752
rect 16568 2737 16632 2752
rect 16632 2737 16648 2752
rect 16648 2737 16712 2752
rect 16712 2737 16728 2752
rect 16728 2737 16758 2752
rect 17182 7648 17418 7710
rect 17182 7584 17212 7648
rect 17212 7584 17228 7648
rect 17228 7584 17292 7648
rect 17292 7584 17308 7648
rect 17308 7584 17372 7648
rect 17372 7584 17388 7648
rect 17388 7584 17418 7648
rect 17182 7474 17418 7584
rect 17182 6115 17418 6351
rect 17182 4756 17418 4992
rect 17182 3397 17418 3633
<< metal5 >>
rect 1056 7710 18908 7752
rect 1056 7474 3865 7710
rect 4101 7474 8304 7710
rect 8540 7474 12743 7710
rect 12979 7474 17182 7710
rect 17418 7474 18908 7710
rect 1056 7432 18908 7474
rect 1056 7050 18908 7092
rect 1056 6814 3205 7050
rect 3441 6814 7644 7050
rect 7880 6814 12083 7050
rect 12319 6814 16522 7050
rect 16758 6814 18908 7050
rect 1056 6772 18908 6814
rect 1056 6351 18908 6393
rect 1056 6115 3865 6351
rect 4101 6115 8304 6351
rect 8540 6115 12743 6351
rect 12979 6115 17182 6351
rect 17418 6115 18908 6351
rect 1056 6073 18908 6115
rect 1056 5691 18908 5733
rect 1056 5455 3205 5691
rect 3441 5455 7644 5691
rect 7880 5455 12083 5691
rect 12319 5455 16522 5691
rect 16758 5455 18908 5691
rect 1056 5413 18908 5455
rect 1056 4992 18908 5034
rect 1056 4756 3865 4992
rect 4101 4756 8304 4992
rect 8540 4756 12743 4992
rect 12979 4756 17182 4992
rect 17418 4756 18908 4992
rect 1056 4714 18908 4756
rect 1056 4332 18908 4374
rect 1056 4096 3205 4332
rect 3441 4096 7644 4332
rect 7880 4096 12083 4332
rect 12319 4096 16522 4332
rect 16758 4096 18908 4332
rect 1056 4054 18908 4096
rect 1056 3633 18908 3675
rect 1056 3397 3865 3633
rect 4101 3397 8304 3633
rect 8540 3397 12743 3633
rect 12979 3397 17182 3633
rect 17418 3397 18908 3633
rect 1056 3355 18908 3397
rect 1056 2973 18908 3015
rect 1056 2737 3205 2973
rect 3441 2737 7644 2973
rect 7880 2737 12083 2973
rect 12319 2737 16522 2973
rect 16758 2737 18908 2973
rect 1056 2695 18908 2737
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 5060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1666464484
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_45
timestamp 1666464484
transform 1 0 5244 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1666464484
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1666464484
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1666464484
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1666464484
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 1666464484
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1666464484
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1666464484
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_70
timestamp 1666464484
transform 1 0 7544 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_78
timestamp 1666464484
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1666464484
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1666464484
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1666464484
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_23
timestamp 1666464484
transform 1 0 3220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_29
timestamp 1666464484
transform 1 0 3772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1666464484
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1666464484
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1666464484
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1666464484
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1666464484
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1666464484
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1666464484
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_99
timestamp 1666464484
transform 1 0 10212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_118
timestamp 1666464484
transform 1 0 11960 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_130
timestamp 1666464484
transform 1 0 13064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_142
timestamp 1666464484
transform 1 0 14168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1666464484
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1666464484
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1666464484
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1666464484
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_43
timestamp 1666464484
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1666464484
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1666464484
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1666464484
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_94
timestamp 1666464484
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1666464484
transform 1 0 10120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_122
timestamp 1666464484
transform 1 0 12328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1666464484
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1666464484
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_22
timestamp 1666464484
transform 1 0 3128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1666464484
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1666464484
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_42
timestamp 1666464484
transform 1 0 4968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1666464484
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1666464484
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_73
timestamp 1666464484
transform 1 0 7820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_79
timestamp 1666464484
transform 1 0 8372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1666464484
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_90
timestamp 1666464484
transform 1 0 9384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_94
timestamp 1666464484
transform 1 0 9752 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_98
timestamp 1666464484
transform 1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1666464484
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_122
timestamp 1666464484
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_129
timestamp 1666464484
transform 1 0 12972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_136
timestamp 1666464484
transform 1 0 13616 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_144
timestamp 1666464484
transform 1 0 14352 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_150
timestamp 1666464484
transform 1 0 14904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_157
timestamp 1666464484
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1666464484
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1666464484
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1666464484
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1666464484
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp 1666464484
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_61
timestamp 1666464484
transform 1 0 6716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1666464484
transform 1 0 7268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1666464484
transform 1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1666464484
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1666464484
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_106
timestamp 1666464484
transform 1 0 10856 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1666464484
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1666464484
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1666464484
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_160
timestamp 1666464484
transform 1 0 15824 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_172
timestamp 1666464484
transform 1 0 16928 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_184
timestamp 1666464484
transform 1 0 18032 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1666464484
transform 1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1666464484
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1666464484
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1666464484
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1666464484
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1666464484
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_61
timestamp 1666464484
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_65
timestamp 1666464484
transform 1 0 7084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_74
timestamp 1666464484
transform 1 0 7912 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_80
timestamp 1666464484
transform 1 0 8464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_84
timestamp 1666464484
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_91
timestamp 1666464484
transform 1 0 9476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1666464484
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_121
timestamp 1666464484
transform 1 0 12236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1666464484
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1666464484
transform 1 0 14444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_152
timestamp 1666464484
transform 1 0 15088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_159
timestamp 1666464484
transform 1 0 15732 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_174
timestamp 1666464484
transform 1 0 17112 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1666464484
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1666464484
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1666464484
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1666464484
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1666464484
transform 1 0 4600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_45
timestamp 1666464484
transform 1 0 5244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1666464484
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 1666464484
transform 1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1666464484
transform 1 0 7268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_74
timestamp 1666464484
transform 1 0 7912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1666464484
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_89
timestamp 1666464484
transform 1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_96
timestamp 1666464484
transform 1 0 9936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_103
timestamp 1666464484
transform 1 0 10580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_110
timestamp 1666464484
transform 1 0 11224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_117
timestamp 1666464484
transform 1 0 11868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_124
timestamp 1666464484
transform 1 0 12512 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1666464484
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1666464484
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1666464484
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp 1666464484
transform 1 0 15824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_167
timestamp 1666464484
transform 1 0 16468 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_174
timestamp 1666464484
transform 1 0 17112 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_181
timestamp 1666464484
transform 1 0 17756 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1666464484
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1666464484
transform 1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1666464484
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_29
timestamp 1666464484
transform 1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_35
timestamp 1666464484
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1666464484
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1666464484
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_70
timestamp 1666464484
transform 1 0 7544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_82
timestamp 1666464484
transform 1 0 8648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1666464484
transform 1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_91
timestamp 1666464484
transform 1 0 9476 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1666464484
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1666464484
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1666464484
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1666464484
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_132
timestamp 1666464484
transform 1 0 13248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1666464484
transform 1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_146
timestamp 1666464484
transform 1 0 14536 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1666464484
transform 1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1666464484
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1666464484
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1666464484
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1666464484
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1666464484
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1666464484
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _029_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _030_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5244 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _031_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _032_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _033_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1666464484
transform -1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _035_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1666464484
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _038_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4140 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _039_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1666464484
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _041_
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _043_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5428 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1666464484
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _045_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7176 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _046_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _047_
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1666464484
transform -1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1666464484
transform -1 0 13616 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp 1666464484
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _051_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7360 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp 1666464484
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _053_
timestamp 1666464484
transform 1 0 11684 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp 1666464484
transform -1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1666464484
transform -1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1666464484
transform -1 0 11960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1666464484
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1666464484
transform -1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _060_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13800 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _061_
timestamp 1666464484
transform 1 0 5612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _062_
timestamp 1666464484
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _063_
timestamp 1666464484
transform 1 0 9108 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _064_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1656 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _065_
timestamp 1666464484
transform 1 0 6808 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _066_
timestamp 1666464484
transform 1 0 10488 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _067_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11224 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _068_
timestamp 1666464484
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6072 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform -1 0 8648 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform -1 0 8648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_9
timestamp 1666464484
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_10
timestamp 1666464484
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_11
timestamp 1666464484
transform -1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_12
timestamp 1666464484
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_13
timestamp 1666464484
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_14
timestamp 1666464484
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_15
timestamp 1666464484
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_16
timestamp 1666464484
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_17
timestamp 1666464484
transform 1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_18
timestamp 1666464484
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_19
timestamp 1666464484
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_20
timestamp 1666464484
transform 1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_21
timestamp 1666464484
transform 1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_22
timestamp 1666464484
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_23
timestamp 1666464484
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_24
timestamp 1666464484
transform 1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_25
timestamp 1666464484
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_26
timestamp 1666464484
transform -1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_27
timestamp 1666464484
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_28
timestamp 1666464484
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_29
timestamp 1666464484
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_30
timestamp 1666464484
transform -1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_31
timestamp 1666464484
transform -1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_32
timestamp 1666464484
transform -1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_33
timestamp 1666464484
transform -1 0 13248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_34
timestamp 1666464484
transform -1 0 13800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_35
timestamp 1666464484
transform -1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_36
timestamp 1666464484
transform -1 0 14444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_37
timestamp 1666464484
transform -1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_38
timestamp 1666464484
transform -1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_39
timestamp 1666464484
transform -1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_40
timestamp 1666464484
transform -1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_41
timestamp 1666464484
transform -1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_42
timestamp 1666464484
transform -1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_43
timestamp 1666464484
transform -1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_44
timestamp 1666464484
transform -1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_45
timestamp 1666464484
transform -1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_46
timestamp 1666464484
transform -1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_47
timestamp 1666464484
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_48
timestamp 1666464484
transform 1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_49
timestamp 1666464484
transform 1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_50
timestamp 1666464484
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_51
timestamp 1666464484
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_52
timestamp 1666464484
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_53
timestamp 1666464484
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_54
timestamp 1666464484
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_55
timestamp 1666464484
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_56
timestamp 1666464484
transform 1 0 8464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_57
timestamp 1666464484
transform -1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_58
timestamp 1666464484
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_59
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_60
timestamp 1666464484
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_61
timestamp 1666464484
transform 1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_62
timestamp 1666464484
transform -1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_63
timestamp 1666464484
transform 1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_64
timestamp 1666464484
transform -1 0 11224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_65
timestamp 1666464484
transform -1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_66
timestamp 1666464484
transform -1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_67
timestamp 1666464484
transform -1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_68
timestamp 1666464484
transform -1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_69
timestamp 1666464484
transform -1 0 14536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_70
timestamp 1666464484
transform -1 0 13800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_71
timestamp 1666464484
transform -1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_72
timestamp 1666464484
transform -1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_73
timestamp 1666464484
transform -1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_74
timestamp 1666464484
transform -1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_75
timestamp 1666464484
transform -1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_76
timestamp 1666464484
transform -1 0 16376 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_77
timestamp 1666464484
transform -1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_78
timestamp 1666464484
transform -1 0 17756 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_wrapper_79
timestamp 1666464484
transform -1 0 15548 0 -1 5440
box -38 -48 314 592
<< labels >>
flabel metal2 s 4710 9200 4766 10000 0 FreeSans 224 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 7470 9200 7526 10000 0 FreeSans 224 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 7746 9200 7802 10000 0 FreeSans 224 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 8022 9200 8078 10000 0 FreeSans 224 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 8298 9200 8354 10000 0 FreeSans 224 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 8574 9200 8630 10000 0 FreeSans 224 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 8850 9200 8906 10000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 9126 9200 9182 10000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 9402 9200 9458 10000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 9678 9200 9734 10000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 9954 9200 10010 10000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 4986 9200 5042 10000 0 FreeSans 224 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 10230 9200 10286 10000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 10506 9200 10562 10000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 10782 9200 10838 10000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 11058 9200 11114 10000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 11334 9200 11390 10000 0 FreeSans 224 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 11610 9200 11666 10000 0 FreeSans 224 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 11886 9200 11942 10000 0 FreeSans 224 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 12162 9200 12218 10000 0 FreeSans 224 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 12438 9200 12494 10000 0 FreeSans 224 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 12714 9200 12770 10000 0 FreeSans 224 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 5262 9200 5318 10000 0 FreeSans 224 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 12990 9200 13046 10000 0 FreeSans 224 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 13266 9200 13322 10000 0 FreeSans 224 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 13542 9200 13598 10000 0 FreeSans 224 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 13818 9200 13874 10000 0 FreeSans 224 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 14094 9200 14150 10000 0 FreeSans 224 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 14370 9200 14426 10000 0 FreeSans 224 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 14646 9200 14702 10000 0 FreeSans 224 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 14922 9200 14978 10000 0 FreeSans 224 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 5538 9200 5594 10000 0 FreeSans 224 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 5814 9200 5870 10000 0 FreeSans 224 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 6090 9200 6146 10000 0 FreeSans 224 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 6366 9200 6422 10000 0 FreeSans 224 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 6642 9200 6698 10000 0 FreeSans 224 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 6918 9200 6974 10000 0 FreeSans 224 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 7194 9200 7250 10000 0 FreeSans 224 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 4802 9200 4858 10000 0 FreeSans 224 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 7562 9200 7618 10000 0 FreeSans 224 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 7838 9200 7894 10000 0 FreeSans 224 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 8114 9200 8170 10000 0 FreeSans 224 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 8390 9200 8446 10000 0 FreeSans 224 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 8666 9200 8722 10000 0 FreeSans 224 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 8942 9200 8998 10000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 9218 9200 9274 10000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 9494 9200 9550 10000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 9770 9200 9826 10000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 10046 9200 10102 10000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 5078 9200 5134 10000 0 FreeSans 224 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 10322 9200 10378 10000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 10598 9200 10654 10000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 10874 9200 10930 10000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11150 9200 11206 10000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 11426 9200 11482 10000 0 FreeSans 224 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 11702 9200 11758 10000 0 FreeSans 224 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 11978 9200 12034 10000 0 FreeSans 224 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 12254 9200 12310 10000 0 FreeSans 224 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 12530 9200 12586 10000 0 FreeSans 224 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 12806 9200 12862 10000 0 FreeSans 224 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 5354 9200 5410 10000 0 FreeSans 224 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 13082 9200 13138 10000 0 FreeSans 224 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 13358 9200 13414 10000 0 FreeSans 224 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 13634 9200 13690 10000 0 FreeSans 224 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 13910 9200 13966 10000 0 FreeSans 224 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 14186 9200 14242 10000 0 FreeSans 224 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 14462 9200 14518 10000 0 FreeSans 224 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 14738 9200 14794 10000 0 FreeSans 224 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 15014 9200 15070 10000 0 FreeSans 224 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 5630 9200 5686 10000 0 FreeSans 224 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 5906 9200 5962 10000 0 FreeSans 224 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 6182 9200 6238 10000 0 FreeSans 224 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 6458 9200 6514 10000 0 FreeSans 224 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 6734 9200 6790 10000 0 FreeSans 224 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 7010 9200 7066 10000 0 FreeSans 224 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 7286 9200 7342 10000 0 FreeSans 224 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4894 9200 4950 10000 0 FreeSans 224 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 7654 9200 7710 10000 0 FreeSans 224 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 7930 9200 7986 10000 0 FreeSans 224 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 8206 9200 8262 10000 0 FreeSans 224 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 8482 9200 8538 10000 0 FreeSans 224 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 8758 9200 8814 10000 0 FreeSans 224 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 9034 9200 9090 10000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 9310 9200 9366 10000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 9586 9200 9642 10000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 9862 9200 9918 10000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 10138 9200 10194 10000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 5170 9200 5226 10000 0 FreeSans 224 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 10414 9200 10470 10000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 10690 9200 10746 10000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 10966 9200 11022 10000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 11242 9200 11298 10000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 11518 9200 11574 10000 0 FreeSans 224 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 11794 9200 11850 10000 0 FreeSans 224 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 12070 9200 12126 10000 0 FreeSans 224 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 12346 9200 12402 10000 0 FreeSans 224 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 12622 9200 12678 10000 0 FreeSans 224 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 12898 9200 12954 10000 0 FreeSans 224 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 5446 9200 5502 10000 0 FreeSans 224 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 13174 9200 13230 10000 0 FreeSans 224 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 13450 9200 13506 10000 0 FreeSans 224 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 13726 9200 13782 10000 0 FreeSans 224 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 14002 9200 14058 10000 0 FreeSans 224 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 14278 9200 14334 10000 0 FreeSans 224 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 14554 9200 14610 10000 0 FreeSans 224 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 14830 9200 14886 10000 0 FreeSans 224 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 15106 9200 15162 10000 0 FreeSans 224 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 5722 9200 5778 10000 0 FreeSans 224 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 5998 9200 6054 10000 0 FreeSans 224 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 6274 9200 6330 10000 0 FreeSans 224 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 6550 9200 6606 10000 0 FreeSans 224 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 6826 9200 6882 10000 0 FreeSans 224 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 7102 9200 7158 10000 0 FreeSans 224 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 7378 9200 7434 10000 0 FreeSans 224 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 3163 2128 3483 7664 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 7602 2128 7922 7664 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 12041 2128 12361 7664 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 16480 2128 16800 7664 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal5 s 1056 2695 18908 3015 0 FreeSans 2560 0 0 0 vccd1
port 114 nsew power bidirectional
flabel metal5 s 1056 4054 18908 4374 0 FreeSans 2560 0 0 0 vccd1
port 114 nsew power bidirectional
flabel metal5 s 1056 5413 18908 5733 0 FreeSans 2560 0 0 0 vccd1
port 114 nsew power bidirectional
flabel metal5 s 1056 6772 18908 7092 0 FreeSans 2560 0 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 3823 2128 4143 7752 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 8262 2128 8582 7752 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 12701 2128 13021 7752 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 17140 2128 17460 7752 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal5 s 1056 3355 18908 3675 0 FreeSans 2560 0 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal5 s 1056 4714 18908 5034 0 FreeSans 2560 0 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal5 s 1056 6073 18908 6393 0 FreeSans 2560 0 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal5 s 1056 7432 18908 7752 0 FreeSans 2560 0 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 9982 7072 9982 7072 0 vccd1
rlabel metal1 9982 7616 9982 7616 0 vssd1
rlabel metal1 9384 4794 9384 4794 0 _000_
rlabel metal1 13202 5338 13202 5338 0 _001_
rlabel metal1 2162 3706 2162 3706 0 _002_
rlabel metal1 6900 3706 6900 3706 0 _003_
rlabel metal1 10810 4488 10810 4488 0 _004_
rlabel metal1 4278 3978 4278 3978 0 _005_
rlabel metal1 5612 5338 5612 5338 0 _006_
rlabel metal1 13662 4794 13662 4794 0 _007_
rlabel metal2 9062 4828 9062 4828 0 _008_
rlabel metal2 3082 4148 3082 4148 0 _009_
rlabel metal1 8602 3706 8602 3706 0 _010_
rlabel metal2 11822 4318 11822 4318 0 _011_
rlabel metal1 12742 4794 12742 4794 0 _012_
rlabel metal1 3036 4114 3036 4114 0 _013_
rlabel metal1 4278 4114 4278 4114 0 _014_
rlabel metal1 7636 5338 7636 5338 0 _015_
rlabel metal2 8878 5134 8878 5134 0 _016_
rlabel metal1 2162 4114 2162 4114 0 _017_
rlabel metal1 5796 4794 5796 4794 0 _018_
rlabel metal1 2530 3536 2530 3536 0 _019_
rlabel metal2 5566 4318 5566 4318 0 _020_
rlabel metal1 5566 3162 5566 3162 0 _021_
rlabel metal1 6164 3502 6164 3502 0 _022_
rlabel metal2 7314 3808 7314 3808 0 _023_
rlabel metal1 7744 3434 7744 3434 0 _024_
rlabel metal1 8372 3638 8372 3638 0 _025_
rlabel metal2 13386 4794 13386 4794 0 _026_
rlabel metal1 9062 4590 9062 4590 0 _027_
rlabel metal1 12581 5202 12581 5202 0 _028_
rlabel metal2 9246 7650 9246 7650 0 io_in[14]
rlabel metal1 5566 4726 5566 4726 0 io_in[5]
rlabel metal1 6210 7378 6210 7378 0 io_in[6]
rlabel metal1 8280 6630 8280 6630 0 io_out[12]
rlabel metal1 8556 7514 8556 7514 0 io_out[13]
rlabel metal1 6992 6630 6992 6630 0 io_out[7]
rlabel metal1 7268 7514 7268 7514 0 io_out[8]
rlabel metal1 1656 4658 1656 4658 0 net1
rlabel metal1 4646 6120 4646 6120 0 net10
rlabel metal2 5750 5066 5750 5066 0 net11
rlabel via2 4370 6851 4370 6851 0 net12
rlabel metal1 2806 6698 2806 6698 0 net13
rlabel metal2 6486 8306 6486 8306 0 net14
rlabel metal1 3956 6766 3956 6766 0 net15
rlabel metal1 4922 7242 4922 7242 0 net16
rlabel metal2 4554 5950 4554 5950 0 net17
rlabel metal1 3450 7412 3450 7412 0 net18
rlabel metal1 6348 6970 6348 6970 0 net19
rlabel metal1 6118 5678 6118 5678 0 net2
rlabel metal1 6118 6766 6118 6766 0 net20
rlabel metal1 7038 6324 7038 6324 0 net21
rlabel metal2 5290 7684 5290 7684 0 net22
rlabel metal1 7084 6834 7084 6834 0 net23
rlabel metal1 8924 5882 8924 5882 0 net24
rlabel metal1 8694 6834 8694 6834 0 net25
rlabel metal1 9844 5202 9844 5202 0 net26
rlabel metal1 9752 6154 9752 6154 0 net27
rlabel metal1 10120 6834 10120 6834 0 net28
rlabel metal1 10580 6834 10580 6834 0 net29
rlabel metal2 12558 4352 12558 4352 0 net3
rlabel metal1 10948 6834 10948 6834 0 net30
rlabel metal1 11454 7378 11454 7378 0 net31
rlabel metal1 11914 7310 11914 7310 0 net32
rlabel metal1 12466 7276 12466 7276 0 net33
rlabel metal1 12995 6766 12995 6766 0 net34
rlabel metal2 12282 8340 12282 8340 0 net35
rlabel metal1 14214 6324 14214 6324 0 net36
rlabel metal1 15272 7242 15272 7242 0 net37
rlabel metal1 14858 6358 14858 6358 0 net38
rlabel metal1 13846 5746 13846 5746 0 net39
rlabel metal2 9982 6290 9982 6290 0 net4
rlabel metal1 14582 6154 14582 6154 0 net40
rlabel metal1 15732 7310 15732 7310 0 net41
rlabel metal1 16836 6902 16836 6902 0 net42
rlabel metal2 18170 7004 18170 7004 0 net43
rlabel metal1 15180 5882 15180 5882 0 net44
rlabel metal1 15962 6290 15962 6290 0 net45
rlabel metal1 4968 3706 4968 3706 0 net46
rlabel metal1 4968 3978 4968 3978 0 net47
rlabel metal1 3680 5202 3680 5202 0 net48
rlabel metal1 2691 6290 2691 6290 0 net49
rlabel metal1 12696 6426 12696 6426 0 net5
rlabel metal1 3634 6086 3634 6086 0 net50
rlabel metal1 6440 4114 6440 4114 0 net51
rlabel metal2 3910 6324 3910 6324 0 net52
rlabel metal1 6762 5236 6762 5236 0 net53
rlabel metal1 5152 6766 5152 6766 0 net54
rlabel metal2 4646 7548 4646 7548 0 net55
rlabel metal1 8740 5202 8740 5202 0 net56
rlabel metal2 9154 6171 9154 6171 0 net57
rlabel metal1 8096 7310 8096 7310 0 net58
rlabel metal1 9200 6290 9200 6290 0 net59
rlabel metal1 6486 6154 6486 6154 0 net6
rlabel metal1 10258 5882 10258 5882 0 net60
rlabel metal1 10120 6290 10120 6290 0 net61
rlabel metal1 10488 6290 10488 6290 0 net62
rlabel metal1 10626 7378 10626 7378 0 net63
rlabel metal2 10994 8340 10994 8340 0 net64
rlabel metal1 11454 6834 11454 6834 0 net65
rlabel metal1 11914 6766 11914 6766 0 net66
rlabel metal2 11822 8068 11822 8068 0 net67
rlabel metal1 12558 7208 12558 7208 0 net68
rlabel metal1 14214 6766 14214 6766 0 net69
rlabel metal2 6670 6630 6670 6630 0 net7
rlabel metal1 13064 5882 13064 5882 0 net70
rlabel metal1 14812 6766 14812 6766 0 net71
rlabel metal1 14444 6970 14444 6970 0 net72
rlabel metal1 15180 6902 15180 6902 0 net73
rlabel metal2 16882 7021 16882 7021 0 net74
rlabel metal1 14490 5814 14490 5814 0 net75
rlabel metal1 15318 6222 15318 6222 0 net76
rlabel metal1 14628 5202 14628 5202 0 net77
rlabel metal1 17526 6732 17526 6732 0 net78
rlabel metal1 15272 5202 15272 5202 0 net79
rlabel metal1 2599 5134 2599 5134 0 net8
rlabel metal1 4094 5066 4094 5066 0 net9
rlabel metal2 11546 5916 11546 5916 0 spi_device.next_state\[0\]
rlabel metal1 2116 3978 2116 3978 0 spi_device.next_state\[1\]
rlabel metal2 13386 5372 13386 5372 0 spi_device.pres_state\[0\]
rlabel metal2 11730 5644 11730 5644 0 spi_device.pres_state\[1\]
rlabel metal1 3956 4522 3956 4522 0 spi_device.t\[0\]
rlabel metal1 5244 4114 5244 4114 0 spi_device.t\[1\]
rlabel metal2 12282 4318 12282 4318 0 spi_device.t\[2\]
<< properties >>
string FIXED_BBOX 0 0 20000 10000
<< end >>
