* NGSPICE file created from spi_register.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_4 abstract view
.subckt sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

.subckt spi_register reg_addr[0] reg_addr[1] reg_addr[2] reg_bus reg_clk reg_data[0]
+ reg_data[1] reg_data[2] reg_data[3] reg_data[4] reg_data[5] reg_data[6] reg_data[7]
+ reg_dir vcc vss
XFILLER_22_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_9_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_66_ reg_bus _03_ vss vss vcc vcc net7 sky130_fd_sc_hd__dlxtn_1
XFILLER_2_132 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_0_57 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_9_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_49_ _15_ _18_ vss vss vcc vcc _23_ sky130_fd_sc_hd__or2_1
XFILLER_18_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
Xoutput7 net7 vss vss vcc vcc reg_data[2] sky130_fd_sc_hd__buf_2
XFILLER_16_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_112 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_3_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_9_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_65_ t\[2\] _15_ vss vss vcc vcc _11_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_2_166 vss vss vcc vcc sky130_fd_sc_hd__fill_2
X_48_ _22_ vss vss vcc vcc _07_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_15_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
Xoutput10 net10 vss vss vcc vcc reg_data[5] sky130_fd_sc_hd__buf_2
Xoutput8 net8 vss vss vcc vcc reg_data[3] sky130_fd_sc_hd__buf_2
XFILLER_16_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_16_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_113 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_69 vss vss vcc vcc sky130_fd_sc_hd__decap_8
X_64_ _13_ _20_ vss vss vcc vcc _10_ sky130_fd_sc_hd__nand2_1
XFILLER_5_120 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_23_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_2_101 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_0_37 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_0_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_145 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_47_ _13_ _18_ vss vss vcc vcc _22_ sky130_fd_sc_hd__or2_1
XFILLER_9_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_1_80 vss vss vcc vcc sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_reg_clk clknet_0_reg_clk vss vss vcc vcc clknet_1_1__leaf_reg_clk sky130_fd_sc_hd__clkbuf_16
Xoutput11 net11 vss vss vcc vcc reg_data[6] sky130_fd_sc_hd__buf_2
Xoutput9 net9 vss vss vcc vcc reg_data[4] sky130_fd_sc_hd__buf_2
XFILLER_16_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XTAP_114 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_90 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_63_ _17_ _27_ _29_ _31_ vss vss vcc vcc _32_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_46_ _21_ vss vss vcc vcc _06_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
Xoutput12 net12 vss vss vcc vcc reg_data[7] sky130_fd_sc_hd__buf_2
XFILLER_15_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_115 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_62_ t\[2\] _30_ vss vss vcc vcc _31_ sky130_fd_sc_hd__and2_1
XFILLER_5_166 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_23_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_125 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_9_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_45_ _18_ _20_ vss vss vcc vcc _21_ sky130_fd_sc_hd__or2_1
XFILLER_6_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_15_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_116 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_81 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_8_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_61_ net9 net10 net11 net12 t\[0\] t\[1\] vss vss vcc vcc _30_ sky130_fd_sc_hd__mux4_1
XFILLER_23_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_82 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_29 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_9_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_44_ t\[1\] t\[0\] vss vss vcc vcc _20_ sky130_fd_sc_hd__or2b_1
XFILLER_1_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_15_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XTAP_106 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_21_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_reg_clk clknet_0_reg_clk vss vss vcc vcc clknet_1_0__leaf_reg_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_8_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_10_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_60_ net7 _13_ _15_ net8 _28_ vss vss vcc vcc _29_ sky130_fd_sc_hd__o221a_1
XFILLER_5_113 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_23_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_94 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_9_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_43_ _19_ vss vss vcc vcc _05_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_1_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_19_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_6_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_107 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_1 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_94 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_23_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_42_ t\[1\] t\[0\] _18_ vss vss vcc vcc _19_ sky130_fd_sc_hd__or3_1
XANTENNA_output5_A net5 vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_18_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_19_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_19_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_108 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_2 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_8_101 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_104 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_4_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_85 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_23_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_118 vss vss vcc vcc sky130_fd_sc_hd__decap_4
X_41_ _17_ _12_ vss vss vcc vcc _18_ sky130_fd_sc_hd__or2_1
XFILLER_20_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_150 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_109 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_22_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XPHY_3 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_16_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_12_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_138 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_2_108 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_4_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_40_ t\[2\] vss vss vcc vcc _17_ sky130_fd_sc_hd__inv_2
XFILLER_13_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_18_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XPHY_4 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_12_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_4_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XANTENNA_input4_A reg_dir vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_24_73 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_1_88 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_1_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_19_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_19_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XANTENNA__59__C net5 vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_10_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_141 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XPHY_5 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_21_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_16_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_137 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_12_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_5_129 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_4_162 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_24_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_6 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_21_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_16_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_141 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_1_166 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_1_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_97 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_1_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_90 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 reg_addr[0] vss vss vcc vcc net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_24_121 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_24_110 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XPHY_7 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_23_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_24_54 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XANTENNA_input2_A reg_addr[1] vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_1_69 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XTAP_91 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 reg_addr[1] vss vss vcc vcc net2 sky130_fd_sc_hd__clkbuf_1
XTAP_80 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_166 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_21_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_16_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_8 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_1_113 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_1_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_92 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 reg_addr[2] vss vss vcc vcc net3 sky130_fd_sc_hd__clkbuf_1
XTAP_70 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_18_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_145 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_15_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_9 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_155 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_13_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_78 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_1_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_93 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 reg_dir vss vss vcc vcc net4 sky130_fd_sc_hd__clkbuf_1
XTAP_60 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_77_ reg_bus _02_ vss vss vcc vcc net6 sky130_fd_sc_hd__dlxtn_1
XTAP_71 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_18_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_113 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_24_102 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_21_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_21_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_131 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_4_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_4_134 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_13_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_92 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_35 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_1_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_76_ clknet_1_1__leaf_reg_clk _11_ vss vss vcc vcc t\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_94 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_83 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_59_ t\[1\] t\[0\] net5 vss vss vcc vcc _28_ sky130_fd_sc_hd__or3_1
XFILLER_21_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_11_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_14_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_1_138 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_1_127 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_1_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_24_69 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_24_47 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_19_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_95 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_75_ clknet_1_0__leaf_reg_clk _10_ vss vss vcc vcc t\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_51 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XTAP_84 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_126 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_58_ net6 _20_ vss vss vcc vcc _27_ sky130_fd_sc_hd__or2_1
XFILLER_21_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_7_144 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_125 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_13_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_96 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_74_ clknet_1_0__leaf_reg_clk _09_ vss vss vcc vcc t\[0\] sky130_fd_sc_hd__dfxtp_2
XTAP_63 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_138 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_21_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_57_ _26_ vss vss vcc vcc _02_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_7_156 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_17_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_5_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XTAP_97 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_73_ reg_bus _01_ vss vss vcc vcc net5 sky130_fd_sc_hd__dlxtn_1
XTAP_53 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_21_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_56_ t\[2\] _12_ _20_ vss vss vcc vcc _26_ sky130_fd_sc_hd__or3_1
XFILLER_23_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_39_ _16_ vss vss vcc vcc _04_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_113 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_17_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_4_116 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_12_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_141 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XTAP_98 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_72_ _32_ _00_ vss vss vcc vcc reg_bus sky130_fd_sc_hd__dlxtn_4
XTAP_65 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_19_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_97 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_2_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_55_ _25_ vss vss vcc vcc _01_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_20_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_20_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_16_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_38_ t\[2\] _12_ _15_ vss vss vcc vcc _16_ sky130_fd_sc_hd__or3_1
XFILLER_22_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_29 vss vss vcc vcc sky130_fd_sc_hd__fill_2
X_71_ reg_bus _08_ vss vss vcc vcc net12 sky130_fd_sc_hd__dlxtn_1
XTAP_99 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_54_ t\[1\] t\[2\] t\[0\] _12_ vss vss vcc vcc _25_ sky130_fd_sc_hd__or4_1
XFILLER_2_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_37_ t\[1\] t\[0\] vss vss vcc vcc _15_ sky130_fd_sc_hd__nand2_1
XFILLER_11_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_97 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_17_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_4_107 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_140 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_14_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_89 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
X_70_ reg_bus _07_ vss vss vcc vcc net11 sky130_fd_sc_hd__dlxtn_1
XTAP_78 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_40 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0_reg_clk_A reg_clk vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_2_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_53_ _24_ vss vss vcc vcc _00_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_36_ _14_ vss vss vcc vcc _03_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_127 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_11_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_8_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_166 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_5_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_5_77 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_10_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_57 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_30 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_52_ net3 net4 net2 net1 vss vss vcc vcc _24_ sky130_fd_sc_hd__or4_1
XFILLER_14_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_35_ t\[2\] _12_ _13_ vss vss vcc vcc _14_ sky130_fd_sc_hd__or3_1
XFILLER_22_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_8_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_0_145 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_14_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_58 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_31 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_20 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_51_ t\[0\] vss vss vcc vcc _09_ sky130_fd_sc_hd__inv_2
XFILLER_23_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_11_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_14_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
X_34_ t\[0\] t\[1\] vss vss vcc vcc _13_ sky130_fd_sc_hd__or2b_1
XFILLER_22_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_3 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_7_107 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_11_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_113 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_90 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_5_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XTAP_59 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XPHY_43 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_18_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_32 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_10 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_21 vss vss vcc vcc sky130_fd_sc_hd__decap_3
X_50_ _23_ vss vss vcc vcc _08_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
X_33_ net3 net2 net1 net4 vss vss vcc vcc _12_ sky130_fd_sc_hd__or4b_2
XFILLER_22_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_11_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_141 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_17_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_3_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_3_166 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_80 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_5_69 vss vss vcc vcc sky130_fd_sc_hd__decap_8
Xclkbuf_0_reg_clk reg_clk vss vss vcc vcc clknet_0_reg_clk sky130_fd_sc_hd__clkbuf_16
XPHY_44 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_33 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_11 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_22 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_2_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_3_91 vss vss vcc vcc sky130_fd_sc_hd__decap_8
XFILLER_11_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_11_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_19_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_164 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_134 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_0_70 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_5_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_12 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_45 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_34 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_2_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_23 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_23_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_6_121 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_8_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_57 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_113 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_124 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_3_146 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_0_138 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_5_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_46 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_35 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_13 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_9_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_24 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_23_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_82 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_8_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_17_69 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_24_3 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_94 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_9_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_47 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_36 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_14 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_25 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_2_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XANTENNA_input3_A reg_addr[2] vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_11_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_112 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_17_15 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_118 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_9_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_48 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_37 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_6_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XPHY_15 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_26 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_11_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_20_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_13_161 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_3_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_22_27 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_0_9 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_6_135 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_8_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_27 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_23_81 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_0_85 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_63 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_0_41 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XPHY_49 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_38 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_27 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_16 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_137 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_15_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_7_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_111 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_10_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_10_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_12_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_17_39 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_117 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_23_93 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_22_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_14_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_6_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_85 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XPHY_17 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_28 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_39 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_17_149 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_17_105 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_22_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_167 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_22_29 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XANTENNA_input1_A reg_addr[0] vss vss vcc vcc sky130_fd_sc_hd__diode_2
XFILLER_10_133 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_3_107 vss vss vcc vcc sky130_fd_sc_hd__decap_4
X_69_ reg_bus _06_ vss vss vcc vcc net10 sky130_fd_sc_hd__dlxtn_1
XFILLER_0_98 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_18_83 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_15_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_29 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XPHY_18 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_15_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_14_109 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_22_153 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_9_113 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_105 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_12_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_68_ reg_bus _05_ vss vss vcc vcc net9 sky130_fd_sc_hd__dlxtn_1
XFILLER_23_51 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_2_141 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_0_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_20_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_65 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XPHY_19 vss vss vcc vcc sky130_fd_sc_hd__decap_3
Xoutput5 net5 vss vss vcc vcc reg_data[0] sky130_fd_sc_hd__buf_2
XTAP_110 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 vss vss vcc vcc sky130_fd_sc_hd__decap_3
XFILLER_22_121 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_3_55 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_3_77 vss vss vcc vcc sky130_fd_sc_hd__fill_2
XFILLER_3_99 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_9_125 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_5_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_128 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_6_139 vss vss vcc vcc sky130_fd_sc_hd__fill_1
XFILLER_12_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_12_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
X_67_ reg_bus _04_ vss vss vcc vcc net8 sky130_fd_sc_hd__dlxtn_1
XFILLER_24_9 vss vss vcc vcc sky130_fd_sc_hd__decap_4
XFILLER_18_85 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_18_41 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_97 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_53 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_20_3 vss vss vcc vcc sky130_ef_sc_hd__decap_12
XFILLER_6_77 vss vss vcc vcc sky130_fd_sc_hd__decap_6
XFILLER_6_99 vss vss vcc vcc sky130_fd_sc_hd__decap_4
Xoutput6 net6 vss vss vcc vcc reg_data[1] sky130_fd_sc_hd__buf_2
XTAP_111 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vss vcc sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vss vss vcc vcc sky130_ef_sc_hd__decap_12
.ends

