VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spi_device
  CLASS BLOCK ;
  FOREIGN spi_device ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN reg_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 246.000 62.930 250.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 246.000 104.330 250.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 246.000 145.730 250.000 ;
    END
  END reg_addr[2]
  PIN reg_bus
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 246.000 187.130 250.000 ;
    END
  END reg_bus
  PIN reg_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 246.000 228.530 250.000 ;
    END
  END reg_clk
  PIN reg_dir
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 246.000 21.530 250.000 ;
    END
  END reg_dir
  PIN spi_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END spi_clk
  PIN spi_miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END spi_miso
  PIN spi_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END spi_mosi
  PIN spi_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END spi_sel
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 5.520 10.640 244.260 236.880 ;
      LAYER met2 ;
        RECT 7.910 245.720 20.970 246.570 ;
        RECT 21.810 245.720 62.370 246.570 ;
        RECT 63.210 245.720 103.770 246.570 ;
        RECT 104.610 245.720 145.170 246.570 ;
        RECT 146.010 245.720 186.570 246.570 ;
        RECT 187.410 245.720 227.970 246.570 ;
        RECT 228.810 245.720 229.900 246.570 ;
        RECT 7.910 10.695 229.900 245.720 ;
      LAYER met3 ;
        RECT 4.000 217.960 176.230 236.805 ;
        RECT 4.400 216.560 176.230 217.960 ;
        RECT 4.000 156.080 176.230 216.560 ;
        RECT 4.400 154.680 176.230 156.080 ;
        RECT 4.000 94.200 176.230 154.680 ;
        RECT 4.400 92.800 176.230 94.200 ;
        RECT 4.000 32.320 176.230 92.800 ;
        RECT 4.400 30.920 176.230 32.320 ;
        RECT 4.000 10.715 176.230 30.920 ;
  END
END spi_device
END LIBRARY

