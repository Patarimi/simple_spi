magic
tech gf180mcuC
magscale 1 10
timestamp 1674139336
<< nwell >>
rect 1258 116384 178726 116902
rect 1258 114816 178726 115680
rect 1258 113248 178726 114112
rect 1258 111680 178726 112544
rect 1258 110112 178726 110976
rect 1258 108544 178726 109408
rect 1258 106976 178726 107840
rect 1258 105408 178726 106272
rect 1258 103840 178726 104704
rect 1258 102272 178726 103136
rect 1258 100704 178726 101568
rect 1258 99136 178726 100000
rect 1258 97568 178726 98432
rect 1258 96000 178726 96864
rect 1258 94432 178726 95296
rect 1258 92864 178726 93728
rect 1258 91296 178726 92160
rect 1258 89728 178726 90592
rect 1258 88160 178726 89024
rect 1258 86592 178726 87456
rect 1258 85024 178726 85888
rect 1258 83456 178726 84320
rect 1258 81888 178726 82752
rect 1258 80320 178726 81184
rect 1258 78752 178726 79616
rect 1258 77184 178726 78048
rect 1258 75616 178726 76480
rect 1258 74048 178726 74912
rect 1258 72480 178726 73344
rect 1258 70912 178726 71776
rect 1258 69344 178726 70208
rect 1258 67776 178726 68640
rect 1258 66208 178726 67072
rect 1258 64640 178726 65504
rect 1258 63072 178726 63936
rect 1258 61504 178726 62368
rect 1258 59936 178726 60800
rect 1258 58368 178726 59232
rect 1258 56800 178726 57664
rect 1258 55232 178726 56096
rect 1258 53664 178726 54528
rect 1258 52096 178726 52960
rect 1258 50528 178726 51392
rect 1258 48960 178726 49824
rect 1258 47392 178726 48256
rect 1258 45824 178726 46688
rect 1258 44256 178726 45120
rect 1258 42688 178726 43552
rect 1258 41120 178726 41984
rect 1258 39552 178726 40416
rect 1258 37984 178726 38848
rect 1258 36416 178726 37280
rect 1258 34848 178726 35712
rect 1258 33280 178726 34144
rect 1258 31712 178726 32576
rect 1258 30144 178726 31008
rect 1258 28576 178726 29440
rect 1258 27008 178726 27872
rect 1258 25440 178726 26304
rect 1258 23872 178726 24736
rect 1258 22304 178726 23168
rect 1258 20736 178726 21600
rect 1258 19168 178726 20032
rect 1258 17600 178726 18464
rect 1258 16032 178726 16896
rect 1258 14464 178726 15328
rect 1258 12896 178726 13760
rect 1258 11353 178726 12192
rect 1258 11328 42680 11353
rect 1258 10599 38717 10624
rect 1258 9785 178726 10599
rect 1258 9760 48168 9785
rect 1258 9031 36632 9056
rect 1258 8217 178726 9031
rect 1258 8192 33608 8217
rect 1258 7463 27560 7488
rect 1258 6649 178726 7463
rect 1258 6624 17928 6649
rect 1258 5895 14568 5920
rect 1258 5081 178726 5895
rect 1258 5056 16429 5081
rect 1258 4327 14680 4352
rect 1258 3513 178726 4327
rect 1258 3488 27224 3513
<< pwell >>
rect 1258 115680 178726 116384
rect 1258 114112 178726 114816
rect 1258 112544 178726 113248
rect 1258 110976 178726 111680
rect 1258 109408 178726 110112
rect 1258 107840 178726 108544
rect 1258 106272 178726 106976
rect 1258 104704 178726 105408
rect 1258 103136 178726 103840
rect 1258 101568 178726 102272
rect 1258 100000 178726 100704
rect 1258 98432 178726 99136
rect 1258 96864 178726 97568
rect 1258 95296 178726 96000
rect 1258 93728 178726 94432
rect 1258 92160 178726 92864
rect 1258 90592 178726 91296
rect 1258 89024 178726 89728
rect 1258 87456 178726 88160
rect 1258 85888 178726 86592
rect 1258 84320 178726 85024
rect 1258 82752 178726 83456
rect 1258 81184 178726 81888
rect 1258 79616 178726 80320
rect 1258 78048 178726 78752
rect 1258 76480 178726 77184
rect 1258 74912 178726 75616
rect 1258 73344 178726 74048
rect 1258 71776 178726 72480
rect 1258 70208 178726 70912
rect 1258 68640 178726 69344
rect 1258 67072 178726 67776
rect 1258 65504 178726 66208
rect 1258 63936 178726 64640
rect 1258 62368 178726 63072
rect 1258 60800 178726 61504
rect 1258 59232 178726 59936
rect 1258 57664 178726 58368
rect 1258 56096 178726 56800
rect 1258 54528 178726 55232
rect 1258 52960 178726 53664
rect 1258 51392 178726 52096
rect 1258 49824 178726 50528
rect 1258 48256 178726 48960
rect 1258 46688 178726 47392
rect 1258 45120 178726 45824
rect 1258 43552 178726 44256
rect 1258 41984 178726 42688
rect 1258 40416 178726 41120
rect 1258 38848 178726 39552
rect 1258 37280 178726 37984
rect 1258 35712 178726 36416
rect 1258 34144 178726 34848
rect 1258 32576 178726 33280
rect 1258 31008 178726 31712
rect 1258 29440 178726 30144
rect 1258 27872 178726 28576
rect 1258 26304 178726 27008
rect 1258 24736 178726 25440
rect 1258 23168 178726 23872
rect 1258 21600 178726 22304
rect 1258 20032 178726 20736
rect 1258 18464 178726 19168
rect 1258 16896 178726 17600
rect 1258 15328 178726 16032
rect 1258 13760 178726 14464
rect 1258 12192 178726 12896
rect 1258 10624 178726 11328
rect 1258 9056 178726 9760
rect 1258 7488 178726 8192
rect 1258 5920 178726 6624
rect 1258 4352 178726 5056
rect 1258 3050 178726 3488
<< obsm1 >>
rect 1344 1710 178640 117570
<< metal2 >>
rect 1344 119200 1456 120000
rect 2912 119200 3024 120000
rect 4480 119200 4592 120000
rect 6048 119200 6160 120000
rect 7616 119200 7728 120000
rect 9184 119200 9296 120000
rect 10752 119200 10864 120000
rect 12320 119200 12432 120000
rect 13888 119200 14000 120000
rect 15456 119200 15568 120000
rect 17024 119200 17136 120000
rect 18592 119200 18704 120000
rect 20160 119200 20272 120000
rect 21728 119200 21840 120000
rect 23296 119200 23408 120000
rect 24864 119200 24976 120000
rect 26432 119200 26544 120000
rect 28000 119200 28112 120000
rect 29568 119200 29680 120000
rect 31136 119200 31248 120000
rect 32704 119200 32816 120000
rect 34272 119200 34384 120000
rect 35840 119200 35952 120000
rect 37408 119200 37520 120000
rect 38976 119200 39088 120000
rect 40544 119200 40656 120000
rect 42112 119200 42224 120000
rect 43680 119200 43792 120000
rect 45248 119200 45360 120000
rect 46816 119200 46928 120000
rect 48384 119200 48496 120000
rect 49952 119200 50064 120000
rect 51520 119200 51632 120000
rect 53088 119200 53200 120000
rect 54656 119200 54768 120000
rect 56224 119200 56336 120000
rect 57792 119200 57904 120000
rect 59360 119200 59472 120000
rect 60928 119200 61040 120000
rect 62496 119200 62608 120000
rect 64064 119200 64176 120000
rect 65632 119200 65744 120000
rect 67200 119200 67312 120000
rect 68768 119200 68880 120000
rect 70336 119200 70448 120000
rect 71904 119200 72016 120000
rect 73472 119200 73584 120000
rect 75040 119200 75152 120000
rect 76608 119200 76720 120000
rect 78176 119200 78288 120000
rect 79744 119200 79856 120000
rect 81312 119200 81424 120000
rect 82880 119200 82992 120000
rect 84448 119200 84560 120000
rect 86016 119200 86128 120000
rect 87584 119200 87696 120000
rect 89152 119200 89264 120000
rect 90720 119200 90832 120000
rect 92288 119200 92400 120000
rect 93856 119200 93968 120000
rect 95424 119200 95536 120000
rect 96992 119200 97104 120000
rect 98560 119200 98672 120000
rect 100128 119200 100240 120000
rect 101696 119200 101808 120000
rect 103264 119200 103376 120000
rect 104832 119200 104944 120000
rect 106400 119200 106512 120000
rect 107968 119200 108080 120000
rect 109536 119200 109648 120000
rect 111104 119200 111216 120000
rect 112672 119200 112784 120000
rect 114240 119200 114352 120000
rect 115808 119200 115920 120000
rect 117376 119200 117488 120000
rect 118944 119200 119056 120000
rect 120512 119200 120624 120000
rect 122080 119200 122192 120000
rect 123648 119200 123760 120000
rect 125216 119200 125328 120000
rect 126784 119200 126896 120000
rect 128352 119200 128464 120000
rect 129920 119200 130032 120000
rect 131488 119200 131600 120000
rect 133056 119200 133168 120000
rect 134624 119200 134736 120000
rect 136192 119200 136304 120000
rect 137760 119200 137872 120000
rect 139328 119200 139440 120000
rect 140896 119200 141008 120000
rect 142464 119200 142576 120000
rect 144032 119200 144144 120000
rect 145600 119200 145712 120000
rect 147168 119200 147280 120000
rect 148736 119200 148848 120000
rect 150304 119200 150416 120000
rect 151872 119200 151984 120000
rect 153440 119200 153552 120000
rect 155008 119200 155120 120000
rect 156576 119200 156688 120000
rect 158144 119200 158256 120000
rect 159712 119200 159824 120000
rect 161280 119200 161392 120000
rect 162848 119200 162960 120000
rect 164416 119200 164528 120000
rect 165984 119200 166096 120000
rect 167552 119200 167664 120000
rect 169120 119200 169232 120000
rect 170688 119200 170800 120000
rect 172256 119200 172368 120000
rect 173824 119200 173936 120000
rect 175392 119200 175504 120000
rect 176960 119200 177072 120000
rect 178528 119200 178640 120000
rect 7280 0 7392 800
rect 7616 0 7728 800
rect 7952 0 8064 800
rect 8288 0 8400 800
rect 8624 0 8736 800
rect 8960 0 9072 800
rect 9296 0 9408 800
rect 9632 0 9744 800
rect 9968 0 10080 800
rect 10304 0 10416 800
rect 10640 0 10752 800
rect 10976 0 11088 800
rect 11312 0 11424 800
rect 11648 0 11760 800
rect 11984 0 12096 800
rect 12320 0 12432 800
rect 12656 0 12768 800
rect 12992 0 13104 800
rect 13328 0 13440 800
rect 13664 0 13776 800
rect 14000 0 14112 800
rect 14336 0 14448 800
rect 14672 0 14784 800
rect 15008 0 15120 800
rect 15344 0 15456 800
rect 15680 0 15792 800
rect 16016 0 16128 800
rect 16352 0 16464 800
rect 16688 0 16800 800
rect 17024 0 17136 800
rect 17360 0 17472 800
rect 17696 0 17808 800
rect 18032 0 18144 800
rect 18368 0 18480 800
rect 18704 0 18816 800
rect 19040 0 19152 800
rect 19376 0 19488 800
rect 19712 0 19824 800
rect 20048 0 20160 800
rect 20384 0 20496 800
rect 20720 0 20832 800
rect 21056 0 21168 800
rect 21392 0 21504 800
rect 21728 0 21840 800
rect 22064 0 22176 800
rect 22400 0 22512 800
rect 22736 0 22848 800
rect 23072 0 23184 800
rect 23408 0 23520 800
rect 23744 0 23856 800
rect 24080 0 24192 800
rect 24416 0 24528 800
rect 24752 0 24864 800
rect 25088 0 25200 800
rect 25424 0 25536 800
rect 25760 0 25872 800
rect 26096 0 26208 800
rect 26432 0 26544 800
rect 26768 0 26880 800
rect 27104 0 27216 800
rect 27440 0 27552 800
rect 27776 0 27888 800
rect 28112 0 28224 800
rect 28448 0 28560 800
rect 28784 0 28896 800
rect 29120 0 29232 800
rect 29456 0 29568 800
rect 29792 0 29904 800
rect 30128 0 30240 800
rect 30464 0 30576 800
rect 30800 0 30912 800
rect 31136 0 31248 800
rect 31472 0 31584 800
rect 31808 0 31920 800
rect 32144 0 32256 800
rect 32480 0 32592 800
rect 32816 0 32928 800
rect 33152 0 33264 800
rect 33488 0 33600 800
rect 33824 0 33936 800
rect 34160 0 34272 800
rect 34496 0 34608 800
rect 34832 0 34944 800
rect 35168 0 35280 800
rect 35504 0 35616 800
rect 35840 0 35952 800
rect 36176 0 36288 800
rect 36512 0 36624 800
rect 36848 0 36960 800
rect 37184 0 37296 800
rect 37520 0 37632 800
rect 37856 0 37968 800
rect 38192 0 38304 800
rect 38528 0 38640 800
rect 38864 0 38976 800
rect 39200 0 39312 800
rect 39536 0 39648 800
rect 39872 0 39984 800
rect 40208 0 40320 800
rect 40544 0 40656 800
rect 40880 0 40992 800
rect 41216 0 41328 800
rect 41552 0 41664 800
rect 41888 0 42000 800
rect 42224 0 42336 800
rect 42560 0 42672 800
rect 42896 0 43008 800
rect 43232 0 43344 800
rect 43568 0 43680 800
rect 43904 0 44016 800
rect 44240 0 44352 800
rect 44576 0 44688 800
rect 44912 0 45024 800
rect 45248 0 45360 800
rect 45584 0 45696 800
rect 45920 0 46032 800
rect 46256 0 46368 800
rect 46592 0 46704 800
rect 46928 0 47040 800
rect 47264 0 47376 800
rect 47600 0 47712 800
rect 47936 0 48048 800
rect 48272 0 48384 800
rect 48608 0 48720 800
rect 48944 0 49056 800
rect 49280 0 49392 800
rect 49616 0 49728 800
rect 49952 0 50064 800
rect 50288 0 50400 800
rect 50624 0 50736 800
rect 50960 0 51072 800
rect 51296 0 51408 800
rect 51632 0 51744 800
rect 51968 0 52080 800
rect 52304 0 52416 800
rect 52640 0 52752 800
rect 52976 0 53088 800
rect 53312 0 53424 800
rect 53648 0 53760 800
rect 53984 0 54096 800
rect 54320 0 54432 800
rect 54656 0 54768 800
rect 54992 0 55104 800
rect 55328 0 55440 800
rect 55664 0 55776 800
rect 56000 0 56112 800
rect 56336 0 56448 800
rect 56672 0 56784 800
rect 57008 0 57120 800
rect 57344 0 57456 800
rect 57680 0 57792 800
rect 58016 0 58128 800
rect 58352 0 58464 800
rect 58688 0 58800 800
rect 59024 0 59136 800
rect 59360 0 59472 800
rect 59696 0 59808 800
rect 60032 0 60144 800
rect 60368 0 60480 800
rect 60704 0 60816 800
rect 61040 0 61152 800
rect 61376 0 61488 800
rect 61712 0 61824 800
rect 62048 0 62160 800
rect 62384 0 62496 800
rect 62720 0 62832 800
rect 63056 0 63168 800
rect 63392 0 63504 800
rect 63728 0 63840 800
rect 64064 0 64176 800
rect 64400 0 64512 800
rect 64736 0 64848 800
rect 65072 0 65184 800
rect 65408 0 65520 800
rect 65744 0 65856 800
rect 66080 0 66192 800
rect 66416 0 66528 800
rect 66752 0 66864 800
rect 67088 0 67200 800
rect 67424 0 67536 800
rect 67760 0 67872 800
rect 68096 0 68208 800
rect 68432 0 68544 800
rect 68768 0 68880 800
rect 69104 0 69216 800
rect 69440 0 69552 800
rect 69776 0 69888 800
rect 70112 0 70224 800
rect 70448 0 70560 800
rect 70784 0 70896 800
rect 71120 0 71232 800
rect 71456 0 71568 800
rect 71792 0 71904 800
rect 72128 0 72240 800
rect 72464 0 72576 800
rect 72800 0 72912 800
rect 73136 0 73248 800
rect 73472 0 73584 800
rect 73808 0 73920 800
rect 74144 0 74256 800
rect 74480 0 74592 800
rect 74816 0 74928 800
rect 75152 0 75264 800
rect 75488 0 75600 800
rect 75824 0 75936 800
rect 76160 0 76272 800
rect 76496 0 76608 800
rect 76832 0 76944 800
rect 77168 0 77280 800
rect 77504 0 77616 800
rect 77840 0 77952 800
rect 78176 0 78288 800
rect 78512 0 78624 800
rect 78848 0 78960 800
rect 79184 0 79296 800
rect 79520 0 79632 800
rect 79856 0 79968 800
rect 80192 0 80304 800
rect 80528 0 80640 800
rect 80864 0 80976 800
rect 81200 0 81312 800
rect 81536 0 81648 800
rect 81872 0 81984 800
rect 82208 0 82320 800
rect 82544 0 82656 800
rect 82880 0 82992 800
rect 83216 0 83328 800
rect 83552 0 83664 800
rect 83888 0 84000 800
rect 84224 0 84336 800
rect 84560 0 84672 800
rect 84896 0 85008 800
rect 85232 0 85344 800
rect 85568 0 85680 800
rect 85904 0 86016 800
rect 86240 0 86352 800
rect 86576 0 86688 800
rect 86912 0 87024 800
rect 87248 0 87360 800
rect 87584 0 87696 800
rect 87920 0 88032 800
rect 88256 0 88368 800
rect 88592 0 88704 800
rect 88928 0 89040 800
rect 89264 0 89376 800
rect 89600 0 89712 800
rect 89936 0 90048 800
rect 90272 0 90384 800
rect 90608 0 90720 800
rect 90944 0 91056 800
rect 91280 0 91392 800
rect 91616 0 91728 800
rect 91952 0 92064 800
rect 92288 0 92400 800
rect 92624 0 92736 800
rect 92960 0 93072 800
rect 93296 0 93408 800
rect 93632 0 93744 800
rect 93968 0 94080 800
rect 94304 0 94416 800
rect 94640 0 94752 800
rect 94976 0 95088 800
rect 95312 0 95424 800
rect 95648 0 95760 800
rect 95984 0 96096 800
rect 96320 0 96432 800
rect 96656 0 96768 800
rect 96992 0 97104 800
rect 97328 0 97440 800
rect 97664 0 97776 800
rect 98000 0 98112 800
rect 98336 0 98448 800
rect 98672 0 98784 800
rect 99008 0 99120 800
rect 99344 0 99456 800
rect 99680 0 99792 800
rect 100016 0 100128 800
rect 100352 0 100464 800
rect 100688 0 100800 800
rect 101024 0 101136 800
rect 101360 0 101472 800
rect 101696 0 101808 800
rect 102032 0 102144 800
rect 102368 0 102480 800
rect 102704 0 102816 800
rect 103040 0 103152 800
rect 103376 0 103488 800
rect 103712 0 103824 800
rect 104048 0 104160 800
rect 104384 0 104496 800
rect 104720 0 104832 800
rect 105056 0 105168 800
rect 105392 0 105504 800
rect 105728 0 105840 800
rect 106064 0 106176 800
rect 106400 0 106512 800
rect 106736 0 106848 800
rect 107072 0 107184 800
rect 107408 0 107520 800
rect 107744 0 107856 800
rect 108080 0 108192 800
rect 108416 0 108528 800
rect 108752 0 108864 800
rect 109088 0 109200 800
rect 109424 0 109536 800
rect 109760 0 109872 800
rect 110096 0 110208 800
rect 110432 0 110544 800
rect 110768 0 110880 800
rect 111104 0 111216 800
rect 111440 0 111552 800
rect 111776 0 111888 800
rect 112112 0 112224 800
rect 112448 0 112560 800
rect 112784 0 112896 800
rect 113120 0 113232 800
rect 113456 0 113568 800
rect 113792 0 113904 800
rect 114128 0 114240 800
rect 114464 0 114576 800
rect 114800 0 114912 800
rect 115136 0 115248 800
rect 115472 0 115584 800
rect 115808 0 115920 800
rect 116144 0 116256 800
rect 116480 0 116592 800
rect 116816 0 116928 800
rect 117152 0 117264 800
rect 117488 0 117600 800
rect 117824 0 117936 800
rect 118160 0 118272 800
rect 118496 0 118608 800
rect 118832 0 118944 800
rect 119168 0 119280 800
rect 119504 0 119616 800
rect 119840 0 119952 800
rect 120176 0 120288 800
rect 120512 0 120624 800
rect 120848 0 120960 800
rect 121184 0 121296 800
rect 121520 0 121632 800
rect 121856 0 121968 800
rect 122192 0 122304 800
rect 122528 0 122640 800
rect 122864 0 122976 800
rect 123200 0 123312 800
rect 123536 0 123648 800
rect 123872 0 123984 800
rect 124208 0 124320 800
rect 124544 0 124656 800
rect 124880 0 124992 800
rect 125216 0 125328 800
rect 125552 0 125664 800
rect 125888 0 126000 800
rect 126224 0 126336 800
rect 126560 0 126672 800
rect 126896 0 127008 800
rect 127232 0 127344 800
rect 127568 0 127680 800
rect 127904 0 128016 800
rect 128240 0 128352 800
rect 128576 0 128688 800
rect 128912 0 129024 800
rect 129248 0 129360 800
rect 129584 0 129696 800
rect 129920 0 130032 800
rect 130256 0 130368 800
rect 130592 0 130704 800
rect 130928 0 131040 800
rect 131264 0 131376 800
rect 131600 0 131712 800
rect 131936 0 132048 800
rect 132272 0 132384 800
rect 132608 0 132720 800
rect 132944 0 133056 800
rect 133280 0 133392 800
rect 133616 0 133728 800
rect 133952 0 134064 800
rect 134288 0 134400 800
rect 134624 0 134736 800
rect 134960 0 135072 800
rect 135296 0 135408 800
rect 135632 0 135744 800
rect 135968 0 136080 800
rect 136304 0 136416 800
rect 136640 0 136752 800
rect 136976 0 137088 800
rect 137312 0 137424 800
rect 137648 0 137760 800
rect 137984 0 138096 800
rect 138320 0 138432 800
rect 138656 0 138768 800
rect 138992 0 139104 800
rect 139328 0 139440 800
rect 139664 0 139776 800
rect 140000 0 140112 800
rect 140336 0 140448 800
rect 140672 0 140784 800
rect 141008 0 141120 800
rect 141344 0 141456 800
rect 141680 0 141792 800
rect 142016 0 142128 800
rect 142352 0 142464 800
rect 142688 0 142800 800
rect 143024 0 143136 800
rect 143360 0 143472 800
rect 143696 0 143808 800
rect 144032 0 144144 800
rect 144368 0 144480 800
rect 144704 0 144816 800
rect 145040 0 145152 800
rect 145376 0 145488 800
rect 145712 0 145824 800
rect 146048 0 146160 800
rect 146384 0 146496 800
rect 146720 0 146832 800
rect 147056 0 147168 800
rect 147392 0 147504 800
rect 147728 0 147840 800
rect 148064 0 148176 800
rect 148400 0 148512 800
rect 148736 0 148848 800
rect 149072 0 149184 800
rect 149408 0 149520 800
rect 149744 0 149856 800
rect 150080 0 150192 800
rect 150416 0 150528 800
rect 150752 0 150864 800
rect 151088 0 151200 800
rect 151424 0 151536 800
rect 151760 0 151872 800
rect 152096 0 152208 800
rect 152432 0 152544 800
rect 152768 0 152880 800
rect 153104 0 153216 800
rect 153440 0 153552 800
rect 153776 0 153888 800
rect 154112 0 154224 800
rect 154448 0 154560 800
rect 154784 0 154896 800
rect 155120 0 155232 800
rect 155456 0 155568 800
rect 155792 0 155904 800
rect 156128 0 156240 800
rect 156464 0 156576 800
rect 156800 0 156912 800
rect 157136 0 157248 800
rect 157472 0 157584 800
rect 157808 0 157920 800
rect 158144 0 158256 800
rect 158480 0 158592 800
rect 158816 0 158928 800
rect 159152 0 159264 800
rect 159488 0 159600 800
rect 159824 0 159936 800
rect 160160 0 160272 800
rect 160496 0 160608 800
rect 160832 0 160944 800
rect 161168 0 161280 800
rect 161504 0 161616 800
rect 161840 0 161952 800
rect 162176 0 162288 800
rect 162512 0 162624 800
rect 162848 0 162960 800
rect 163184 0 163296 800
rect 163520 0 163632 800
rect 163856 0 163968 800
rect 164192 0 164304 800
rect 164528 0 164640 800
rect 164864 0 164976 800
rect 165200 0 165312 800
rect 165536 0 165648 800
rect 165872 0 165984 800
rect 166208 0 166320 800
rect 166544 0 166656 800
rect 166880 0 166992 800
rect 167216 0 167328 800
rect 167552 0 167664 800
rect 167888 0 168000 800
rect 168224 0 168336 800
rect 168560 0 168672 800
rect 168896 0 169008 800
rect 169232 0 169344 800
rect 169568 0 169680 800
rect 169904 0 170016 800
rect 170240 0 170352 800
rect 170576 0 170688 800
rect 170912 0 171024 800
rect 171248 0 171360 800
rect 171584 0 171696 800
rect 171920 0 172032 800
rect 172256 0 172368 800
rect 172592 0 172704 800
<< obsm2 >>
rect 3084 119140 4420 119364
rect 4652 119140 5988 119364
rect 6220 119140 7556 119364
rect 7788 119140 9124 119364
rect 9356 119140 10692 119364
rect 10924 119140 12260 119364
rect 12492 119140 13828 119364
rect 14060 119140 15396 119364
rect 15628 119140 16964 119364
rect 17196 119140 18532 119364
rect 18764 119140 20100 119364
rect 20332 119140 21668 119364
rect 21900 119140 23236 119364
rect 23468 119140 24804 119364
rect 25036 119140 26372 119364
rect 26604 119140 27940 119364
rect 28172 119140 29508 119364
rect 29740 119140 31076 119364
rect 31308 119140 32644 119364
rect 32876 119140 34212 119364
rect 34444 119140 35780 119364
rect 36012 119140 37348 119364
rect 37580 119140 38916 119364
rect 39148 119140 40484 119364
rect 40716 119140 42052 119364
rect 42284 119140 43620 119364
rect 43852 119140 45188 119364
rect 45420 119140 46756 119364
rect 46988 119140 48324 119364
rect 48556 119140 49892 119364
rect 50124 119140 51460 119364
rect 51692 119140 53028 119364
rect 53260 119140 54596 119364
rect 54828 119140 56164 119364
rect 56396 119140 57732 119364
rect 57964 119140 59300 119364
rect 59532 119140 60868 119364
rect 61100 119140 62436 119364
rect 62668 119140 64004 119364
rect 64236 119140 65572 119364
rect 65804 119140 67140 119364
rect 67372 119140 68708 119364
rect 68940 119140 70276 119364
rect 70508 119140 71844 119364
rect 72076 119140 73412 119364
rect 73644 119140 74980 119364
rect 75212 119140 76548 119364
rect 76780 119140 78116 119364
rect 78348 119140 79684 119364
rect 79916 119140 81252 119364
rect 81484 119140 82820 119364
rect 83052 119140 84388 119364
rect 84620 119140 85956 119364
rect 86188 119140 87524 119364
rect 87756 119140 89092 119364
rect 89324 119140 90660 119364
rect 90892 119140 92228 119364
rect 92460 119140 93796 119364
rect 94028 119140 95364 119364
rect 95596 119140 96932 119364
rect 97164 119140 98500 119364
rect 98732 119140 100068 119364
rect 100300 119140 101636 119364
rect 101868 119140 103204 119364
rect 103436 119140 104772 119364
rect 105004 119140 106340 119364
rect 106572 119140 107908 119364
rect 108140 119140 109476 119364
rect 109708 119140 111044 119364
rect 111276 119140 112612 119364
rect 112844 119140 114180 119364
rect 114412 119140 115748 119364
rect 115980 119140 117316 119364
rect 117548 119140 118884 119364
rect 119116 119140 120452 119364
rect 120684 119140 122020 119364
rect 122252 119140 123588 119364
rect 123820 119140 125156 119364
rect 125388 119140 126724 119364
rect 126956 119140 128292 119364
rect 128524 119140 129860 119364
rect 130092 119140 131428 119364
rect 131660 119140 132996 119364
rect 133228 119140 134564 119364
rect 134796 119140 136132 119364
rect 136364 119140 137700 119364
rect 137932 119140 139268 119364
rect 139500 119140 140836 119364
rect 141068 119140 142404 119364
rect 142636 119140 143972 119364
rect 144204 119140 145540 119364
rect 145772 119140 147108 119364
rect 147340 119140 148676 119364
rect 148908 119140 150244 119364
rect 150476 119140 151812 119364
rect 152044 119140 153380 119364
rect 153612 119140 154948 119364
rect 155180 119140 156516 119364
rect 156748 119140 158084 119364
rect 158316 119140 159652 119364
rect 159884 119140 161220 119364
rect 161452 119140 162788 119364
rect 163020 119140 164356 119364
rect 164588 119140 165924 119364
rect 166156 119140 167492 119364
rect 167724 119140 169060 119364
rect 169292 119140 170628 119364
rect 170860 119140 172196 119364
rect 172428 119140 173764 119364
rect 173996 119140 175332 119364
rect 175564 119140 176900 119364
rect 177132 119140 178468 119364
rect 2940 860 178612 119140
rect 2940 800 7220 860
rect 7452 800 7556 860
rect 7788 800 7892 860
rect 8124 800 8228 860
rect 8460 800 8564 860
rect 8796 800 8900 860
rect 9132 800 9236 860
rect 9468 800 9572 860
rect 9804 800 9908 860
rect 10140 800 10244 860
rect 10476 800 10580 860
rect 10812 800 10916 860
rect 11148 800 11252 860
rect 11484 800 11588 860
rect 11820 800 11924 860
rect 12156 800 12260 860
rect 12492 800 12596 860
rect 12828 800 12932 860
rect 13164 800 13268 860
rect 13500 800 13604 860
rect 13836 800 13940 860
rect 14172 800 14276 860
rect 14508 800 14612 860
rect 14844 800 14948 860
rect 15180 800 15284 860
rect 15516 800 15620 860
rect 15852 800 15956 860
rect 16188 800 16292 860
rect 16524 800 16628 860
rect 16860 800 16964 860
rect 17196 800 17300 860
rect 17532 800 17636 860
rect 17868 800 17972 860
rect 18204 800 18308 860
rect 18540 800 18644 860
rect 18876 800 18980 860
rect 19212 800 19316 860
rect 19548 800 19652 860
rect 19884 800 19988 860
rect 20220 800 20324 860
rect 20556 800 20660 860
rect 20892 800 20996 860
rect 21228 800 21332 860
rect 21564 800 21668 860
rect 21900 800 22004 860
rect 22236 800 22340 860
rect 22572 800 22676 860
rect 22908 800 23012 860
rect 23244 800 23348 860
rect 23580 800 23684 860
rect 23916 800 24020 860
rect 24252 800 24356 860
rect 24588 800 24692 860
rect 24924 800 25028 860
rect 25260 800 25364 860
rect 25596 800 25700 860
rect 25932 800 26036 860
rect 26268 800 26372 860
rect 26604 800 26708 860
rect 26940 800 27044 860
rect 27276 800 27380 860
rect 27612 800 27716 860
rect 27948 800 28052 860
rect 28284 800 28388 860
rect 28620 800 28724 860
rect 28956 800 29060 860
rect 29292 800 29396 860
rect 29628 800 29732 860
rect 29964 800 30068 860
rect 30300 800 30404 860
rect 30636 800 30740 860
rect 30972 800 31076 860
rect 31308 800 31412 860
rect 31644 800 31748 860
rect 31980 800 32084 860
rect 32316 800 32420 860
rect 32652 800 32756 860
rect 32988 800 33092 860
rect 33324 800 33428 860
rect 33660 800 33764 860
rect 33996 800 34100 860
rect 34332 800 34436 860
rect 34668 800 34772 860
rect 35004 800 35108 860
rect 35340 800 35444 860
rect 35676 800 35780 860
rect 36012 800 36116 860
rect 36348 800 36452 860
rect 36684 800 36788 860
rect 37020 800 37124 860
rect 37356 800 37460 860
rect 37692 800 37796 860
rect 38028 800 38132 860
rect 38364 800 38468 860
rect 38700 800 38804 860
rect 39036 800 39140 860
rect 39372 800 39476 860
rect 39708 800 39812 860
rect 40044 800 40148 860
rect 40380 800 40484 860
rect 40716 800 40820 860
rect 41052 800 41156 860
rect 41388 800 41492 860
rect 41724 800 41828 860
rect 42060 800 42164 860
rect 42396 800 42500 860
rect 42732 800 42836 860
rect 43068 800 43172 860
rect 43404 800 43508 860
rect 43740 800 43844 860
rect 44076 800 44180 860
rect 44412 800 44516 860
rect 44748 800 44852 860
rect 45084 800 45188 860
rect 45420 800 45524 860
rect 45756 800 45860 860
rect 46092 800 46196 860
rect 46428 800 46532 860
rect 46764 800 46868 860
rect 47100 800 47204 860
rect 47436 800 47540 860
rect 47772 800 47876 860
rect 48108 800 48212 860
rect 48444 800 48548 860
rect 48780 800 48884 860
rect 49116 800 49220 860
rect 49452 800 49556 860
rect 49788 800 49892 860
rect 50124 800 50228 860
rect 50460 800 50564 860
rect 50796 800 50900 860
rect 51132 800 51236 860
rect 51468 800 51572 860
rect 51804 800 51908 860
rect 52140 800 52244 860
rect 52476 800 52580 860
rect 52812 800 52916 860
rect 53148 800 53252 860
rect 53484 800 53588 860
rect 53820 800 53924 860
rect 54156 800 54260 860
rect 54492 800 54596 860
rect 54828 800 54932 860
rect 55164 800 55268 860
rect 55500 800 55604 860
rect 55836 800 55940 860
rect 56172 800 56276 860
rect 56508 800 56612 860
rect 56844 800 56948 860
rect 57180 800 57284 860
rect 57516 800 57620 860
rect 57852 800 57956 860
rect 58188 800 58292 860
rect 58524 800 58628 860
rect 58860 800 58964 860
rect 59196 800 59300 860
rect 59532 800 59636 860
rect 59868 800 59972 860
rect 60204 800 60308 860
rect 60540 800 60644 860
rect 60876 800 60980 860
rect 61212 800 61316 860
rect 61548 800 61652 860
rect 61884 800 61988 860
rect 62220 800 62324 860
rect 62556 800 62660 860
rect 62892 800 62996 860
rect 63228 800 63332 860
rect 63564 800 63668 860
rect 63900 800 64004 860
rect 64236 800 64340 860
rect 64572 800 64676 860
rect 64908 800 65012 860
rect 65244 800 65348 860
rect 65580 800 65684 860
rect 65916 800 66020 860
rect 66252 800 66356 860
rect 66588 800 66692 860
rect 66924 800 67028 860
rect 67260 800 67364 860
rect 67596 800 67700 860
rect 67932 800 68036 860
rect 68268 800 68372 860
rect 68604 800 68708 860
rect 68940 800 69044 860
rect 69276 800 69380 860
rect 69612 800 69716 860
rect 69948 800 70052 860
rect 70284 800 70388 860
rect 70620 800 70724 860
rect 70956 800 71060 860
rect 71292 800 71396 860
rect 71628 800 71732 860
rect 71964 800 72068 860
rect 72300 800 72404 860
rect 72636 800 72740 860
rect 72972 800 73076 860
rect 73308 800 73412 860
rect 73644 800 73748 860
rect 73980 800 74084 860
rect 74316 800 74420 860
rect 74652 800 74756 860
rect 74988 800 75092 860
rect 75324 800 75428 860
rect 75660 800 75764 860
rect 75996 800 76100 860
rect 76332 800 76436 860
rect 76668 800 76772 860
rect 77004 800 77108 860
rect 77340 800 77444 860
rect 77676 800 77780 860
rect 78012 800 78116 860
rect 78348 800 78452 860
rect 78684 800 78788 860
rect 79020 800 79124 860
rect 79356 800 79460 860
rect 79692 800 79796 860
rect 80028 800 80132 860
rect 80364 800 80468 860
rect 80700 800 80804 860
rect 81036 800 81140 860
rect 81372 800 81476 860
rect 81708 800 81812 860
rect 82044 800 82148 860
rect 82380 800 82484 860
rect 82716 800 82820 860
rect 83052 800 83156 860
rect 83388 800 83492 860
rect 83724 800 83828 860
rect 84060 800 84164 860
rect 84396 800 84500 860
rect 84732 800 84836 860
rect 85068 800 85172 860
rect 85404 800 85508 860
rect 85740 800 85844 860
rect 86076 800 86180 860
rect 86412 800 86516 860
rect 86748 800 86852 860
rect 87084 800 87188 860
rect 87420 800 87524 860
rect 87756 800 87860 860
rect 88092 800 88196 860
rect 88428 800 88532 860
rect 88764 800 88868 860
rect 89100 800 89204 860
rect 89436 800 89540 860
rect 89772 800 89876 860
rect 90108 800 90212 860
rect 90444 800 90548 860
rect 90780 800 90884 860
rect 91116 800 91220 860
rect 91452 800 91556 860
rect 91788 800 91892 860
rect 92124 800 92228 860
rect 92460 800 92564 860
rect 92796 800 92900 860
rect 93132 800 93236 860
rect 93468 800 93572 860
rect 93804 800 93908 860
rect 94140 800 94244 860
rect 94476 800 94580 860
rect 94812 800 94916 860
rect 95148 800 95252 860
rect 95484 800 95588 860
rect 95820 800 95924 860
rect 96156 800 96260 860
rect 96492 800 96596 860
rect 96828 800 96932 860
rect 97164 800 97268 860
rect 97500 800 97604 860
rect 97836 800 97940 860
rect 98172 800 98276 860
rect 98508 800 98612 860
rect 98844 800 98948 860
rect 99180 800 99284 860
rect 99516 800 99620 860
rect 99852 800 99956 860
rect 100188 800 100292 860
rect 100524 800 100628 860
rect 100860 800 100964 860
rect 101196 800 101300 860
rect 101532 800 101636 860
rect 101868 800 101972 860
rect 102204 800 102308 860
rect 102540 800 102644 860
rect 102876 800 102980 860
rect 103212 800 103316 860
rect 103548 800 103652 860
rect 103884 800 103988 860
rect 104220 800 104324 860
rect 104556 800 104660 860
rect 104892 800 104996 860
rect 105228 800 105332 860
rect 105564 800 105668 860
rect 105900 800 106004 860
rect 106236 800 106340 860
rect 106572 800 106676 860
rect 106908 800 107012 860
rect 107244 800 107348 860
rect 107580 800 107684 860
rect 107916 800 108020 860
rect 108252 800 108356 860
rect 108588 800 108692 860
rect 108924 800 109028 860
rect 109260 800 109364 860
rect 109596 800 109700 860
rect 109932 800 110036 860
rect 110268 800 110372 860
rect 110604 800 110708 860
rect 110940 800 111044 860
rect 111276 800 111380 860
rect 111612 800 111716 860
rect 111948 800 112052 860
rect 112284 800 112388 860
rect 112620 800 112724 860
rect 112956 800 113060 860
rect 113292 800 113396 860
rect 113628 800 113732 860
rect 113964 800 114068 860
rect 114300 800 114404 860
rect 114636 800 114740 860
rect 114972 800 115076 860
rect 115308 800 115412 860
rect 115644 800 115748 860
rect 115980 800 116084 860
rect 116316 800 116420 860
rect 116652 800 116756 860
rect 116988 800 117092 860
rect 117324 800 117428 860
rect 117660 800 117764 860
rect 117996 800 118100 860
rect 118332 800 118436 860
rect 118668 800 118772 860
rect 119004 800 119108 860
rect 119340 800 119444 860
rect 119676 800 119780 860
rect 120012 800 120116 860
rect 120348 800 120452 860
rect 120684 800 120788 860
rect 121020 800 121124 860
rect 121356 800 121460 860
rect 121692 800 121796 860
rect 122028 800 122132 860
rect 122364 800 122468 860
rect 122700 800 122804 860
rect 123036 800 123140 860
rect 123372 800 123476 860
rect 123708 800 123812 860
rect 124044 800 124148 860
rect 124380 800 124484 860
rect 124716 800 124820 860
rect 125052 800 125156 860
rect 125388 800 125492 860
rect 125724 800 125828 860
rect 126060 800 126164 860
rect 126396 800 126500 860
rect 126732 800 126836 860
rect 127068 800 127172 860
rect 127404 800 127508 860
rect 127740 800 127844 860
rect 128076 800 128180 860
rect 128412 800 128516 860
rect 128748 800 128852 860
rect 129084 800 129188 860
rect 129420 800 129524 860
rect 129756 800 129860 860
rect 130092 800 130196 860
rect 130428 800 130532 860
rect 130764 800 130868 860
rect 131100 800 131204 860
rect 131436 800 131540 860
rect 131772 800 131876 860
rect 132108 800 132212 860
rect 132444 800 132548 860
rect 132780 800 132884 860
rect 133116 800 133220 860
rect 133452 800 133556 860
rect 133788 800 133892 860
rect 134124 800 134228 860
rect 134460 800 134564 860
rect 134796 800 134900 860
rect 135132 800 135236 860
rect 135468 800 135572 860
rect 135804 800 135908 860
rect 136140 800 136244 860
rect 136476 800 136580 860
rect 136812 800 136916 860
rect 137148 800 137252 860
rect 137484 800 137588 860
rect 137820 800 137924 860
rect 138156 800 138260 860
rect 138492 800 138596 860
rect 138828 800 138932 860
rect 139164 800 139268 860
rect 139500 800 139604 860
rect 139836 800 139940 860
rect 140172 800 140276 860
rect 140508 800 140612 860
rect 140844 800 140948 860
rect 141180 800 141284 860
rect 141516 800 141620 860
rect 141852 800 141956 860
rect 142188 800 142292 860
rect 142524 800 142628 860
rect 142860 800 142964 860
rect 143196 800 143300 860
rect 143532 800 143636 860
rect 143868 800 143972 860
rect 144204 800 144308 860
rect 144540 800 144644 860
rect 144876 800 144980 860
rect 145212 800 145316 860
rect 145548 800 145652 860
rect 145884 800 145988 860
rect 146220 800 146324 860
rect 146556 800 146660 860
rect 146892 800 146996 860
rect 147228 800 147332 860
rect 147564 800 147668 860
rect 147900 800 148004 860
rect 148236 800 148340 860
rect 148572 800 148676 860
rect 148908 800 149012 860
rect 149244 800 149348 860
rect 149580 800 149684 860
rect 149916 800 150020 860
rect 150252 800 150356 860
rect 150588 800 150692 860
rect 150924 800 151028 860
rect 151260 800 151364 860
rect 151596 800 151700 860
rect 151932 800 152036 860
rect 152268 800 152372 860
rect 152604 800 152708 860
rect 152940 800 153044 860
rect 153276 800 153380 860
rect 153612 800 153716 860
rect 153948 800 154052 860
rect 154284 800 154388 860
rect 154620 800 154724 860
rect 154956 800 155060 860
rect 155292 800 155396 860
rect 155628 800 155732 860
rect 155964 800 156068 860
rect 156300 800 156404 860
rect 156636 800 156740 860
rect 156972 800 157076 860
rect 157308 800 157412 860
rect 157644 800 157748 860
rect 157980 800 158084 860
rect 158316 800 158420 860
rect 158652 800 158756 860
rect 158988 800 159092 860
rect 159324 800 159428 860
rect 159660 800 159764 860
rect 159996 800 160100 860
rect 160332 800 160436 860
rect 160668 800 160772 860
rect 161004 800 161108 860
rect 161340 800 161444 860
rect 161676 800 161780 860
rect 162012 800 162116 860
rect 162348 800 162452 860
rect 162684 800 162788 860
rect 163020 800 163124 860
rect 163356 800 163460 860
rect 163692 800 163796 860
rect 164028 800 164132 860
rect 164364 800 164468 860
rect 164700 800 164804 860
rect 165036 800 165140 860
rect 165372 800 165476 860
rect 165708 800 165812 860
rect 166044 800 166148 860
rect 166380 800 166484 860
rect 166716 800 166820 860
rect 167052 800 167156 860
rect 167388 800 167492 860
rect 167724 800 167828 860
rect 168060 800 168164 860
rect 168396 800 168500 860
rect 168732 800 168836 860
rect 169068 800 169172 860
rect 169404 800 169508 860
rect 169740 800 169844 860
rect 170076 800 170180 860
rect 170412 800 170516 860
rect 170748 800 170852 860
rect 171084 800 171188 860
rect 171420 800 171524 860
rect 171756 800 171860 860
rect 172092 800 172196 860
rect 172428 800 172532 860
rect 172764 800 178612 860
<< obsm3 >>
rect 2930 28 173710 117572
<< metal4 >>
rect 4448 3076 4768 116876
rect 19808 3076 20128 116876
rect 35168 3076 35488 116876
rect 50528 3076 50848 116876
rect 65888 3076 66208 116876
rect 81248 3076 81568 116876
rect 96608 3076 96928 116876
rect 111968 3076 112288 116876
rect 127328 3076 127648 116876
rect 142688 3076 143008 116876
rect 158048 3076 158368 116876
rect 173408 3076 173728 116876
<< obsm4 >>
rect 23100 3016 35108 116238
rect 35548 3016 50468 116238
rect 50908 3016 65828 116238
rect 66268 3016 81188 116238
rect 81628 3016 96548 116238
rect 96988 3016 111908 116238
rect 112348 3016 114548 116238
rect 23100 18 114548 3016
<< labels >>
rlabel metal2 s 1344 119200 1456 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 48384 119200 48496 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 53088 119200 53200 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57792 119200 57904 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 62496 119200 62608 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 67200 119200 67312 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71904 119200 72016 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 76608 119200 76720 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81312 119200 81424 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86016 119200 86128 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 90720 119200 90832 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6048 119200 6160 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95424 119200 95536 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100128 119200 100240 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104832 119200 104944 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 109536 119200 109648 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114240 119200 114352 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118944 119200 119056 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 123648 119200 123760 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 128352 119200 128464 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 133056 119200 133168 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 137760 119200 137872 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10752 119200 10864 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 142464 119200 142576 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 147168 119200 147280 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 151872 119200 151984 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 156576 119200 156688 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 161280 119200 161392 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 165984 119200 166096 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 170688 119200 170800 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 175392 119200 175504 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 15456 119200 15568 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 20160 119200 20272 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24864 119200 24976 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29568 119200 29680 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 34272 119200 34384 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38976 119200 39088 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 43680 119200 43792 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2912 119200 3024 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 49952 119200 50064 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 54656 119200 54768 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 59360 119200 59472 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 64064 119200 64176 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68768 119200 68880 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 73472 119200 73584 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 78176 119200 78288 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82880 119200 82992 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 87584 119200 87696 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92288 119200 92400 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7616 119200 7728 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 96992 119200 97104 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 101696 119200 101808 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 106400 119200 106512 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 111104 119200 111216 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 115808 119200 115920 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 120512 119200 120624 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 125216 119200 125328 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 129920 119200 130032 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 134624 119200 134736 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 139328 119200 139440 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12320 119200 12432 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 144032 119200 144144 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 148736 119200 148848 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 153440 119200 153552 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 158144 119200 158256 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 162848 119200 162960 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 167552 119200 167664 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 172256 119200 172368 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 176960 119200 177072 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 17024 119200 17136 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21728 119200 21840 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 26432 119200 26544 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 31136 119200 31248 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35840 119200 35952 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 40544 119200 40656 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 45248 119200 45360 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4480 119200 4592 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 51520 119200 51632 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 56224 119200 56336 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 60928 119200 61040 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 65632 119200 65744 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 70336 119200 70448 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 75040 119200 75152 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 79744 119200 79856 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 84448 119200 84560 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 89152 119200 89264 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93856 119200 93968 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9184 119200 9296 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 98560 119200 98672 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 103264 119200 103376 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 107968 119200 108080 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 112672 119200 112784 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 117376 119200 117488 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 122080 119200 122192 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 126784 119200 126896 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 131488 119200 131600 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 136192 119200 136304 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 140896 119200 141008 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13888 119200 14000 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 145600 119200 145712 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 150304 119200 150416 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 155008 119200 155120 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 159712 119200 159824 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 164416 119200 164528 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 169120 119200 169232 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 173824 119200 173936 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 178528 119200 178640 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18592 119200 18704 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 23296 119200 23408 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 28000 119200 28112 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32704 119200 32816 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37408 119200 37520 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 42112 119200 42224 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46816 119200 46928 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 171920 0 172032 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 172256 0 172368 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 172592 0 172704 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 42896 0 43008 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 143696 0 143808 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 144704 0 144816 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 145712 0 145824 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 146720 0 146832 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 147728 0 147840 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 148736 0 148848 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 149744 0 149856 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 150752 0 150864 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 151760 0 151872 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 152768 0 152880 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 52976 0 53088 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 153776 0 153888 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 154784 0 154896 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 155792 0 155904 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 156800 0 156912 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 157808 0 157920 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 158816 0 158928 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 159824 0 159936 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 160832 0 160944 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 161840 0 161952 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 162848 0 162960 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 53984 0 54096 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 163856 0 163968 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 164864 0 164976 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 165872 0 165984 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 166880 0 166992 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 167888 0 168000 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 168896 0 169008 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 169904 0 170016 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 170912 0 171024 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 54992 0 55104 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 56000 0 56112 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 57008 0 57120 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 58016 0 58128 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 59024 0 59136 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 60032 0 60144 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 61040 0 61152 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 62048 0 62160 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 43904 0 44016 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 63056 0 63168 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 64064 0 64176 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 65072 0 65184 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 66080 0 66192 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 67088 0 67200 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 68096 0 68208 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 69104 0 69216 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 70112 0 70224 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 71120 0 71232 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 72128 0 72240 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 44912 0 45024 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 73136 0 73248 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 74144 0 74256 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 75152 0 75264 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 76160 0 76272 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 77168 0 77280 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 78176 0 78288 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 79184 0 79296 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 80192 0 80304 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 81200 0 81312 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 82208 0 82320 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 45920 0 46032 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 83216 0 83328 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 84224 0 84336 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 85232 0 85344 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86240 0 86352 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87248 0 87360 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88256 0 88368 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89264 0 89376 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90272 0 90384 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91280 0 91392 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 92288 0 92400 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 46928 0 47040 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 93296 0 93408 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 94304 0 94416 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 95312 0 95424 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 96320 0 96432 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 97328 0 97440 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 98336 0 98448 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 99344 0 99456 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 100352 0 100464 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 101360 0 101472 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 102368 0 102480 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 47936 0 48048 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 103376 0 103488 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 104384 0 104496 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 105392 0 105504 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 106400 0 106512 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 107408 0 107520 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 108416 0 108528 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 109424 0 109536 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 110432 0 110544 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 111440 0 111552 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 112448 0 112560 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 48944 0 49056 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 113456 0 113568 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 114464 0 114576 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 115472 0 115584 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 116480 0 116592 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 117488 0 117600 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 118496 0 118608 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 119504 0 119616 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 120512 0 120624 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 121520 0 121632 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 122528 0 122640 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 49952 0 50064 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 123536 0 123648 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 124544 0 124656 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 125552 0 125664 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 126560 0 126672 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 127568 0 127680 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 128576 0 128688 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 129584 0 129696 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 130592 0 130704 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 131600 0 131712 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 132608 0 132720 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 50960 0 51072 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 133616 0 133728 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 134624 0 134736 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 135632 0 135744 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 136640 0 136752 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 137648 0 137760 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 138656 0 138768 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 139664 0 139776 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 140672 0 140784 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 141680 0 141792 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 142688 0 142800 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 51968 0 52080 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 43232 0 43344 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 144032 0 144144 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 145040 0 145152 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 146048 0 146160 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 147056 0 147168 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 148064 0 148176 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 149072 0 149184 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 150080 0 150192 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 151088 0 151200 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 152096 0 152208 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 153104 0 153216 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 53312 0 53424 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 154112 0 154224 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 155120 0 155232 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 156128 0 156240 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 157136 0 157248 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 158144 0 158256 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 159152 0 159264 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 160160 0 160272 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 161168 0 161280 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 162176 0 162288 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 163184 0 163296 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 54320 0 54432 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 164192 0 164304 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 165200 0 165312 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 166208 0 166320 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 167216 0 167328 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 168224 0 168336 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 169232 0 169344 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 170240 0 170352 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 171248 0 171360 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 55328 0 55440 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 56336 0 56448 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 57344 0 57456 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 58352 0 58464 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 59360 0 59472 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 60368 0 60480 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 61376 0 61488 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 62384 0 62496 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 44240 0 44352 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 63392 0 63504 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 64400 0 64512 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 65408 0 65520 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 66416 0 66528 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 67424 0 67536 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 68432 0 68544 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 69440 0 69552 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 70448 0 70560 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 71456 0 71568 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 72464 0 72576 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 45248 0 45360 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 73472 0 73584 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 74480 0 74592 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 75488 0 75600 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 76496 0 76608 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 77504 0 77616 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 78512 0 78624 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 79520 0 79632 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 80528 0 80640 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 81536 0 81648 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 82544 0 82656 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 46256 0 46368 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 83552 0 83664 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 84560 0 84672 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 85568 0 85680 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 86576 0 86688 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 87584 0 87696 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88592 0 88704 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 89600 0 89712 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 90608 0 90720 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 91616 0 91728 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 92624 0 92736 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 47264 0 47376 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 93632 0 93744 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 94640 0 94752 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 95648 0 95760 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 96656 0 96768 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 97664 0 97776 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 98672 0 98784 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 99680 0 99792 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 100688 0 100800 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 101696 0 101808 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 102704 0 102816 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 48272 0 48384 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 103712 0 103824 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 104720 0 104832 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 105728 0 105840 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 106736 0 106848 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 107744 0 107856 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 108752 0 108864 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 109760 0 109872 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 110768 0 110880 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 111776 0 111888 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 112784 0 112896 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 49280 0 49392 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 113792 0 113904 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 114800 0 114912 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 115808 0 115920 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 116816 0 116928 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 117824 0 117936 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 118832 0 118944 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 119840 0 119952 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 120848 0 120960 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 121856 0 121968 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 122864 0 122976 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 50288 0 50400 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 123872 0 123984 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 124880 0 124992 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 125888 0 126000 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 126896 0 127008 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 127904 0 128016 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 128912 0 129024 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 129920 0 130032 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 130928 0 131040 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 131936 0 132048 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 132944 0 133056 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 51296 0 51408 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 133952 0 134064 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 134960 0 135072 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 135968 0 136080 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 136976 0 137088 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 137984 0 138096 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 138992 0 139104 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 140000 0 140112 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 141008 0 141120 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 142016 0 142128 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 143024 0 143136 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 52304 0 52416 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 43568 0 43680 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 144368 0 144480 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 145376 0 145488 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 146384 0 146496 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 147392 0 147504 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 148400 0 148512 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 149408 0 149520 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 150416 0 150528 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 151424 0 151536 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 152432 0 152544 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 153440 0 153552 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 53648 0 53760 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 154448 0 154560 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 155456 0 155568 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 156464 0 156576 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 157472 0 157584 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 158480 0 158592 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 159488 0 159600 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 160496 0 160608 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 161504 0 161616 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 162512 0 162624 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 163520 0 163632 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 54656 0 54768 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 164528 0 164640 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 165536 0 165648 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 166544 0 166656 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 167552 0 167664 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 168560 0 168672 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 169568 0 169680 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 170576 0 170688 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 171584 0 171696 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 55664 0 55776 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 56672 0 56784 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 57680 0 57792 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 58688 0 58800 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 59696 0 59808 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 60704 0 60816 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 61712 0 61824 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 62720 0 62832 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 44576 0 44688 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 63728 0 63840 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 64736 0 64848 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 65744 0 65856 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 66752 0 66864 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 67760 0 67872 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 68768 0 68880 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 69776 0 69888 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 70784 0 70896 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 71792 0 71904 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 72800 0 72912 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 45584 0 45696 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 73808 0 73920 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 74816 0 74928 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 75824 0 75936 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 76832 0 76944 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 77840 0 77952 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 78848 0 78960 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 79856 0 79968 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80864 0 80976 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 81872 0 81984 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 82880 0 82992 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 46592 0 46704 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 83888 0 84000 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 84896 0 85008 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 85904 0 86016 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 86912 0 87024 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 87920 0 88032 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 88928 0 89040 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 89936 0 90048 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 90944 0 91056 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 91952 0 92064 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 92960 0 93072 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 47600 0 47712 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 93968 0 94080 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 94976 0 95088 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 95984 0 96096 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 96992 0 97104 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 98000 0 98112 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 99008 0 99120 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 100016 0 100128 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 101024 0 101136 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 102032 0 102144 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 103040 0 103152 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 48608 0 48720 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 104048 0 104160 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 105056 0 105168 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 106064 0 106176 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 107072 0 107184 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 108080 0 108192 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 109088 0 109200 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 110096 0 110208 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 111104 0 111216 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 112112 0 112224 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 113120 0 113232 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 49616 0 49728 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 114128 0 114240 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 115136 0 115248 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 116144 0 116256 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 117152 0 117264 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 118160 0 118272 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 119168 0 119280 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 120176 0 120288 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 121184 0 121296 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 122192 0 122304 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 123200 0 123312 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 50624 0 50736 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 124208 0 124320 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 125216 0 125328 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 126224 0 126336 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 127232 0 127344 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 128240 0 128352 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 129248 0 129360 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 130256 0 130368 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 131264 0 131376 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 132272 0 132384 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 133280 0 133392 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 51632 0 51744 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 134288 0 134400 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 135296 0 135408 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 136304 0 136416 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 137312 0 137424 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 138320 0 138432 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 139328 0 139440 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 140336 0 140448 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 141344 0 141456 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 142352 0 142464 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 143360 0 143472 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 52640 0 52752 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4448 3076 4768 116876 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 116876 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 116876 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 116876 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 116876 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 116876 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 116876 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 116876 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 116876 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 116876 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 116876 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 116876 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 7280 0 7392 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 7616 0 7728 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 7952 0 8064 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 9296 0 9408 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 20720 0 20832 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 21728 0 21840 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 22736 0 22848 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 23744 0 23856 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 24752 0 24864 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 25760 0 25872 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 26768 0 26880 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 27776 0 27888 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 28784 0 28896 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 29792 0 29904 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 10640 0 10752 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 30800 0 30912 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 31808 0 31920 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 32816 0 32928 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 33824 0 33936 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 34832 0 34944 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 35840 0 35952 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 36848 0 36960 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 37856 0 37968 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 38864 0 38976 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 39872 0 39984 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 11984 0 12096 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 40880 0 40992 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 41888 0 42000 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 13328 0 13440 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 14672 0 14784 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 15680 0 15792 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 16688 0 16800 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 17696 0 17808 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 18704 0 18816 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 19712 0 19824 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 8288 0 8400 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 9632 0 9744 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 21056 0 21168 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 22064 0 22176 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 23072 0 23184 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 24080 0 24192 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 25088 0 25200 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 26096 0 26208 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 27104 0 27216 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 28112 0 28224 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 29120 0 29232 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 30128 0 30240 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 10976 0 11088 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 31136 0 31248 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 32144 0 32256 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 33152 0 33264 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 34160 0 34272 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 35168 0 35280 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 36176 0 36288 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 37184 0 37296 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 38192 0 38304 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 39200 0 39312 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 40208 0 40320 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 12320 0 12432 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 41216 0 41328 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 42224 0 42336 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 13664 0 13776 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 15008 0 15120 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 16016 0 16128 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 17024 0 17136 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 18032 0 18144 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 19040 0 19152 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 20048 0 20160 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 9968 0 10080 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 21392 0 21504 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 22400 0 22512 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 23408 0 23520 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 24416 0 24528 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 25424 0 25536 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 26432 0 26544 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 27440 0 27552 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 28448 0 28560 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 29456 0 29568 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 30464 0 30576 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 11312 0 11424 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 31472 0 31584 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 32480 0 32592 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 33488 0 33600 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 34496 0 34608 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 35504 0 35616 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 36512 0 36624 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 37520 0 37632 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 38528 0 38640 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 39536 0 39648 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 40544 0 40656 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 12656 0 12768 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 41552 0 41664 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 42560 0 42672 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 14000 0 14112 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 15344 0 15456 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 16352 0 16464 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 17360 0 17472 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 18368 0 18480 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 19376 0 19488 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 20384 0 20496 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 10304 0 10416 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 11648 0 11760 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 12992 0 13104 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 14336 0 14448 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 8624 0 8736 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 8960 0 9072 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3903776
string GDS_FILE /home/mpotereau/DigitalFlowTest/gf_spi_test/openlane/user_proj_example/runs/23_01_19_15_39/results/signoff/user_proj_example.magic.gds
string GDS_START 264624
<< end >>

