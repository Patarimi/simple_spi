magic
tech sky130A
magscale 1 2
timestamp 1680689121
<< nwell >>
rect 1066 20933 22854 21499
rect 1066 19845 22854 20411
rect 1066 18757 22854 19323
rect 1066 17669 22854 18235
rect 1066 16581 22854 17147
rect 1066 15493 22854 16059
rect 1066 14405 22854 14971
rect 1066 13317 22854 13883
rect 1066 12229 22854 12795
rect 1066 11141 22854 11707
rect 1066 10053 22854 10619
rect 1066 8965 22854 9531
rect 1066 7877 22854 8443
rect 1066 6789 22854 7355
rect 1066 5701 22854 6267
rect 1066 4613 22854 5179
rect 1066 3525 22854 4091
rect 1066 2437 22854 3003
<< obsli1 >>
rect 1104 2159 22816 21777
<< obsm1 >>
rect 1104 2128 22976 21808
<< metal2 >>
rect 1674 23200 1730 24000
rect 4618 23200 4674 24000
rect 7562 23200 7618 24000
rect 10506 23200 10562 24000
rect 13450 23200 13506 24000
rect 16394 23200 16450 24000
rect 19338 23200 19394 24000
rect 22282 23200 22338 24000
rect 2042 0 2098 800
rect 5998 0 6054 800
rect 9954 0 10010 800
rect 13910 0 13966 800
rect 17866 0 17922 800
rect 21822 0 21878 800
<< obsm2 >>
rect 1786 23144 4562 23338
rect 4730 23144 7506 23338
rect 7674 23144 10450 23338
rect 10618 23144 13394 23338
rect 13562 23144 16338 23338
rect 16506 23144 19282 23338
rect 19450 23144 22226 23338
rect 22394 23144 22970 23338
rect 1730 856 22970 23144
rect 1730 800 1986 856
rect 2154 800 5942 856
rect 6110 800 9898 856
rect 10066 800 13854 856
rect 14022 800 17810 856
rect 17978 800 21766 856
rect 21934 800 22970 856
<< obsm3 >>
rect 3660 2143 22974 21793
<< metal4 >>
rect 3658 2128 3978 21808
rect 6372 2128 6692 21808
rect 9086 2128 9406 21808
rect 11800 2128 12120 21808
rect 14514 2128 14834 21808
rect 17228 2128 17548 21808
rect 19942 2128 20262 21808
rect 22656 2128 22976 21808
<< labels >>
rlabel metal2 s 5998 0 6054 800 6 reg_addr[0]
port 1 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 reg_addr[1]
port 2 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 reg_addr[2]
port 3 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 reg_bus
port 4 nsew signal bidirectional
rlabel metal2 s 21822 0 21878 800 6 reg_clk
port 5 nsew signal input
rlabel metal2 s 1674 23200 1730 24000 6 reg_data[0]
port 6 nsew signal output
rlabel metal2 s 4618 23200 4674 24000 6 reg_data[1]
port 7 nsew signal output
rlabel metal2 s 7562 23200 7618 24000 6 reg_data[2]
port 8 nsew signal output
rlabel metal2 s 10506 23200 10562 24000 6 reg_data[3]
port 9 nsew signal output
rlabel metal2 s 13450 23200 13506 24000 6 reg_data[4]
port 10 nsew signal output
rlabel metal2 s 16394 23200 16450 24000 6 reg_data[5]
port 11 nsew signal output
rlabel metal2 s 19338 23200 19394 24000 6 reg_data[6]
port 12 nsew signal output
rlabel metal2 s 22282 23200 22338 24000 6 reg_data[7]
port 13 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 reg_dir
port 14 nsew signal input
rlabel metal4 s 3658 2128 3978 21808 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 9086 2128 9406 21808 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 14514 2128 14834 21808 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 19942 2128 20262 21808 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 6372 2128 6692 21808 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 11800 2128 12120 21808 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 17228 2128 17548 21808 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 22656 2128 22976 21808 6 vssd1
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 563730
string GDS_FILE /home/mpotereau/DigitalFlowTest/ol_mpw2304c/openlane/spi_register/runs/23_04_05_12_03/results/signoff/spi_register.magic.gds
string GDS_START 201088
<< end >>

