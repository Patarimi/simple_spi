magic
tech sky130A
magscale 1 2
timestamp 1673535537
<< obsli1 >>
rect 1104 2159 16836 15793
<< obsm1 >>
rect 1104 2128 16995 15824
<< metal2 >>
rect 1582 17200 1638 18000
rect 4526 17200 4582 18000
rect 7470 17200 7526 18000
rect 10414 17200 10470 18000
rect 13358 17200 13414 18000
rect 16302 17200 16358 18000
<< obsm2 >>
rect 1490 17144 1526 17354
rect 1694 17144 4470 17354
rect 4638 17144 7414 17354
rect 7582 17144 10358 17354
rect 10526 17144 13302 17354
rect 13470 17144 16246 17354
rect 16414 17144 16989 17354
rect 1490 2139 16989 17144
<< metal3 >>
rect 0 15648 800 15768
rect 0 11160 800 11280
rect 0 6672 800 6792
rect 0 2184 800 2304
<< obsm3 >>
rect 880 15568 16993 15809
rect 800 11360 16993 15568
rect 880 11080 16993 11360
rect 800 6872 16993 11080
rect 880 6592 16993 6872
rect 800 2384 16993 6592
rect 880 2143 16993 2384
<< metal4 >>
rect 2910 2128 3230 15824
rect 4876 2128 5196 15824
rect 6843 2128 7163 15824
rect 8809 2128 9129 15824
rect 10776 2128 11096 15824
rect 12742 2128 13062 15824
rect 14709 2128 15029 15824
rect 16675 2128 16995 15824
<< labels >>
rlabel metal2 s 4526 17200 4582 18000 6 reg_addr[0]
port 1 nsew signal output
rlabel metal2 s 7470 17200 7526 18000 6 reg_addr[1]
port 2 nsew signal output
rlabel metal2 s 10414 17200 10470 18000 6 reg_addr[2]
port 3 nsew signal output
rlabel metal2 s 13358 17200 13414 18000 6 reg_bus
port 4 nsew signal bidirectional
rlabel metal2 s 16302 17200 16358 18000 6 reg_clk
port 5 nsew signal output
rlabel metal2 s 1582 17200 1638 18000 6 reg_dir
port 6 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 spi_clk
port 7 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 spi_miso
port 8 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 spi_mosi
port 9 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 spi_sel
port 10 nsew signal input
rlabel metal4 s 2910 2128 3230 15824 6 vcc
port 11 nsew power bidirectional
rlabel metal4 s 6843 2128 7163 15824 6 vcc
port 11 nsew power bidirectional
rlabel metal4 s 10776 2128 11096 15824 6 vcc
port 11 nsew power bidirectional
rlabel metal4 s 14709 2128 15029 15824 6 vcc
port 11 nsew power bidirectional
rlabel metal4 s 4876 2128 5196 15824 6 vss
port 12 nsew ground bidirectional
rlabel metal4 s 8809 2128 9129 15824 6 vss
port 12 nsew ground bidirectional
rlabel metal4 s 12742 2128 13062 15824 6 vss
port 12 nsew ground bidirectional
rlabel metal4 s 16675 2128 16995 15824 6 vss
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 463486
string GDS_FILE /home/mpotereau/DigitalFlowTest/gf_spi_test/openlane/spi_device/runs/23_01_12_15_57/results/signoff/spi_device.magic.gds
string GDS_START 205272
<< end >>

